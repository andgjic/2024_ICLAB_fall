/**************************************************************************/
// Copyright (c) 2024, OASIS Lab
// MODULE: PATTERN
// FILE NAME: PATTERN.v
// VERSRION: 1.0
// DATE: August 15, 2024
// AUTHOR: Yu-Hsuan Hsu, NYCU IEE
// DESCRIPTION: ICLAB2024FALL / LAB3 / PATTERN
// MODIFICATION HISTORY:
// Date                 Description
// 
/**************************************************************************/

`ifdef RTL
    `define CYCLE_TIME 40.0
`endif
`ifdef GATE
    `define CYCLE_TIME 40.0
`endif

module PATTERN(
	//OUTPUT
	rst_n,
	clk,
	in_valid,
	tetrominoes,
	position,
	//INPUT
	tetris_valid,
	score_valid,
	fail,
	score,
	tetris
);


`protected
>eE<U?4]A;]A,Hb<22dL#Q-<[g\YcbbV3\[.M6(3>GGD]>\D?)?Y,)]9ULf5?0P9
eC=_e[XENH>VUZO+:Yb72L:f9DEC+[51If.GcW@P2PDf>fCQP0,1_H&[I3R(89]d
R3Y+be1C0Ob[,gX?/<VEd337IOMgAVN-C6]V#\B4E5.RK.8ATA>J&]aV8ATFJG&a
<1+b5<Pg#gYKV?&H)DW6EFJe@66]WfZBT._VB;_P^;)-cCCM6(BDSD[QeD:\SaI/
V>F&/L5J6L^/7Df<ZLR<>H<)_(.V8D>&([LR/HXO_1[^47e^Pe2OS;[QK$
`endprotected
output reg			rst_n, clk, in_valid;
output reg	[2:0]	tetrominoes;
output reg  [2:0]	position;
input 				tetris_valid, score_valid, fail;
input 		[3:0]	score;
input		[71:0]	tetris;


`protected
a,Jc2KK73>1ZR)JYc3(+0I2._O+B=g=8W8#5dE(]7V41f;NNde31&)IZ.=TZb@4c
^5f]g..M;(LdJ\R.WV;V^gZK5W:GI&&M_E#CTM/FDCI+^&;AZUBG4#O_Ec]L?M&M
#XR8)_@7U54UJ7ObV2RPa[6<A_e_\;W-Lf1)S1FeRMWER[W7EEb>AZ+63cF3^Z#:
d])-;+dXVBPf#)G)badD?&Y_-35bc?H[3I11?0aIX-A@FOAE6B+N)2T=b:6W.0g6
9N0K(]5,TfffNV=Y;6Z[S>^;GGOZ(0@g)XP?>QESNL@@?U.T/+/V,=OdaY&VR#Q+
F7;f4)R9g=A1<9Hc&f8CKbK0g04S=g](&d[/+S[I4/?>f+c54\5bI9_1J^\c3CC+
[g[D,BSddDPSe9832OTSJI?.gVN=2:&\0D<WH4N_F5X<b<3&[(MO3+OR:-SN^0bO
bT>?C0;:U4IeNLLRO5GCWU1Qcd23E8JL+E3+>SE?&#+=f9V7M6_IdG=#QGXL51C1
1PQEd=AJ#&2#O7.S:Y.E?.9EU7V(.Eb9(b+3/9:6X5aUNT:9K0:K/dCW\eW6]NJK
IQd:#\L0?=2(1Y;Q]Q)YQ8.<CQ82LG3D^dfQAgMT:__-^/(2@AL[2#9IDWX0F;6M
W1?,?/Zg&afLCL^L-]0M<QRc6ZeYgG-U3DJf+1#He<e^Af9P#4f4.L0(T4XOBgC.
FLI_MWLE?#7f6XXH3PA;^_Yg60Z(ONdL2_Ub1R;CZcO6[)R7(;Qa.ggTWOg1BceN
_-,F2)\WdRS09TdX/ZI\M^d(#&Me2/1M+PF#0>cN#@E,EK_/K7^,Y;-&Z+>cHbbZ
REg]?\g9XB?R.fL&VS&TO(TJL;LEQ)V2^2;QgTR.U:)8AO2&aQ[+[091H]#_YH5,
ZdFf_RF#9GRG6[.DOLeJL10I(e4LI1OM-_e2HeEP?PaAfJJ0J3KP/8HDT=/C)65@
LBVf5UM/9;eQOW].BR+WRDfPb90XUFcA:RKA0RL,3&;a0I_cB5WZ;>1_A-0aK-IC
;53SQJQ+=L@,gYbA3M^+8F/3-9d(A;GDAZ_@gVM1D>3MT#W=01TD6T/V.<e5WfDA
7L2d/Q_Q>Q[)U2/HXR7&]=-4WNeBWMdD+D-3^K>f<[cc-4S++OC2R9;C<8(G#LKT
<H5,PNU.SS903NCee&b&&[4GFU.#REOUL91\GaU7@/MJ3SY?ScB^d92HZ5fMM\2I
AZb#,5Z3?ZQ>2CB\[YO<8affZd,KKOFgD:b9E\c)5A/)MT978UJV,/=?:VaeGVG&
;:KMOY3<B334[5:\_M?Lc/<9,F-W3,^+0dFV-ZQ6)?9:H)_.8=\Z?J[^&/8&C3?^
(48^SdK6=#.&F5aPJZS..W53J,SP3)PWV1[J>R8f?d?M]CA^@2V8/\(?)4Ba#00A
S/)CKHTNP;+]&QIAQ6/>.\NdK\.U]UR7R6e7<51.-PffBLE]a\/6B_]42L6D8#,f
1S9L(KWOKA/e^c_Mg:LWEQ+()MgbI9cP_;J6K:O<Ya8D0=fD[T.aXa-,&UQ6P)DD
/3VEHbX@TC;/[;&VHa#4D58H^P__+)Z:94>d=_7.WF7M9=YOF2BJU/IGBEL,I;=e
^E1X^J.Y=]c6HU^R\-_-ZZA3/U/CSB[e,D/&3.+1#7I-e#:X\XNd<HR1:NI]HI&F
E=TYa?//F-N4T.(Z?]7+.6B/<VKRXd^L]EO<3[gK/:O_SM6c_1+=DAEUR#f+1>d.
1aKH^X)-3Y/5ZWWX>^QUMZLQ98DQb@+X(XF\&aA)K&)R96_8^-/0F-66[C1T1=5,
RMOg4e[Q_MWf4E=\K(.d>NC,2bC\f>0>efN11^UQWE[))S]D=I0-3(7.[#H3E4,P
]>6EY41/L-4UB2-Z#fM2_YKd(F5PQGKDL-.V68A08cg=9X?fB+>\bIUO[#WA=H9F
a4X>+-4;6I5B1#-g-HB^54La3?H7d0_LeE)#>71eB<V\.\^fMC?gH_6#\FOf>b[,
_.=U0X[EB#9U19J6J:N:B9R05116.=5>.LO]?6CR<&F1dEdD;1b5H;c2,1Saf3[R
<REQXJ9E,\,,5Cf(A=)X2:<(_F7<8P[)(R.QbRV<Db-E#^O6dfV,c2;Qa4Jb(0\D
;J)VYV1W<SUBe4>a//5?.?J>C9A.OZJ/KY:gJBdGYZTCaBNb2gT&K/J<^S<(P>E9
g:SF(I#WPC,Mb6dR\M51ZG-R4>Dc(_\3b)(_]G1OEGL;9?1MN]cK?:5g/5368PIW
WVO7B5gAd6?Jg)bB-[^VTZGABK:W1R1bW2Ca-]D,)(;MYSN>PbG?L7c2LQ0^X4+\
Y6GeY&^9DZa+J4HL.2>7;[^]Ab679JTKFVOWG/I?,ce:8B/,5GD3NU4bSDJT,V5U
@BE3Cg&/V:--#B&>^Z7HR00fJ4R(TN8PZR>+]+I9[IWA9.)BHFQdGS.0MPdI;97V
W8E2&QMS2e/g^J1BTL6QMI?S_53A82(4]&H=X#AQ\]Pdcg4[?I_SO7A\d_\]K-[1
.1&e63^;g/A+X_YVVM+N(KLI,fE#0R91S?EWS?aFO#6fEBb3.&MY^&bZc4A1b[CI
E/d4[3c?B[B[<1)Za,Wc&KQ8.NRP5P@bDZa&Nc<^WG<-H]BC[&Y,(^2N@ZJ0CL17
5I8dKZ:ATU;GH^1b<F73;#AR@)a_0A?<#Zde2HQJ?Z]G?Yf?VH+^N)6>S/IC&OWE
[fb>f>:H,1(.g8_81X):=YaI,,4M^54])eT3>94)S,acM40X/1f[1?3=629?_RX@
E<>FFbJ](0^D[0>V]?UI-+GSVcO4WZ7eeTdfJ0+2_1d2K5?M^+=DJeOK^33QR1D2
&5fNX>LGcOC1+>F3TddC;)b@ba,K1P&N0Q&/1KGC-8\3;ENd1aa=a\5)VXaVA[EO
(ZJZSR?B&<B:-7Nf+GZ=)CAS)_TYc#a10:?:(MYe/-/K^8,)[F,A4=Xb(f)LT^N:
MP[TB06TH[:NfOOX0(7SLL<UNg^+_6>ffHSLa?&G>eIMeA+DHYRM<80ND&1#T8Gb
b/JE6/S2I<T^3(13M@T;EOU\?:G)?^,T_)RI=@I#PO;>Y?[BQ8.FdYeGI\+;P81<
))VZ_+8985=e?\8^;I:gF;2b:0L1:5J#6a_6d_e+G[;>E]MUbc#F+a-JISB?.WdF
Q?:@dZ^QY8FWEU-)f,0:R?g]C>Od@J?4)b5D6_DU=\YQGGdWGG;ISGW3LCfAS)+I
9T#4?:bcC,N3ZT69e@^PSH#W_GDF_;WVNZZTLH7ScL<X=@=00IF[QCLT,1dg4&O.
?-R?:9B=AVSFY<I.NA&<]Xd-^L2.S/?^\B2#GNS5XK4S,.IRWYO/]ae[3?\aYQO#
-2f>KWHL<B_]REf?,R>:)I[@KcSSL/@),N0UHPOcgK9&b@=b,c,Sg1F[5.NbO-OW
_M>;_KNHa+;N/5g6A4\BV5c[B0-]EY?fR)]\b?cVE[2SMS,-CcgBd1WHYO^\1+RP
C:g\Y2Z7[e>OU1dTaK>1==DJF(+,6Y)9PB#W9T&=SD#D+4.R+7>+&<eCZZ5GS>?;
Q(QS>WdMPd_Hf]?0DL<]S#Ng:#4P&DI1>F,=aLQB+4:#5V,IG=;@RAW3PIKC-LIN
_C(LS+YdFJaHJD8FKO>:8GO:_J;Qc,Na@)P8U,a0)3&c03<GRZ-2#Q3V+4ITHTIb
D)HJG-gB=Q6L.&34[DQ.]GP0)2-9^GgZ8e\M,PA3Ufd7TL9gA5f<Q@Y&2I?J;[M6
f4DT^(16O9QG8IFK4Gc-\\T09R_XL,DG0U&56MWPE2RLN5S2@f@701XU1KeUM(OA
:?8IVBS]Be6[A\9[;4>X1AR\SdN&G,RVCQ>@66&CR##V@[M?L(7_Z,ENDL:Y7gU:
/9#4SOHb^>1VY45_&OIQ1(31_f3#56E7G;4ab4/-KJ:,NPQCL+8AFM0H7Af3@:be
aBSK)+T^HJg^ON#HJ#Y:MONDE;G#L?Sa_#B6F;R>dCK+]T+)()BCf5Q;7]CN4a@;
1S14cQ;92.T8(W6[6?=JQJ+DYYSdT;ZT<6d=Q9#ZbSF;(1EKL?T]87,MSNI/=>:P
_&0X:N,)<1G<5<_?L#b=O0]DAB-]8&TC=&ffK+NMJ?gaN;M>,gW6FE;IPaVRA/<V
XUT&^0G&GcY/S;Bgd68L.C:@+0KPQHa\6/F#-9e)(=<_a&S]B&J7\>(aM-Fg2(8e
<JU5cG&CbG(>e+1_g70^5DK=C.W.c0KZUabeGO6C4^B0N:NMMZ96;_C:>XLHc5I.
TRgIEE0#S(?X\T,Z[D^SYN@)ET.VdO(/#&@4>L]6&:/#Z:OJSe2/=QcUe8e<,-03
.]J5HM=++^:AMDb6?cQfU:UNWB4B2BP0KRPA6[IR:#F.?Ada1MP9#P[aR_6=82-a
BA>=&XVK^#O,^g)\?FGG]#f__<G@\QKSVPOAMKV:R[9SW>R6N-3b:J5S&9+J.8(-
SQZZ46XFHeF3g/&<a<X55eFQ4;RA+/cR/4QH]Mb?QD2[Y/A]0SJ6d3BNU587cX??
U2G+3O(UGR.]9Q/fe,^W>(M^V+baQCSW.,]#&GRC+(ZVS_ZW)=C;@BM]@Y=ZJb7/
M@JIZ?Q4TZg:#[]ZYCb6-@bOLM.9Z1Q;6cQdFCfJ[.CE1cJfF=G_K/::U\[5-G:M
2C#M\Z9P(N>\=-aA./?#/ZYC=dD>7DWN3N6TO=(U-WZ88IGD0f-f04C_?UcbB/#Y
cOEGY93gIF9ATG&FcXRfd+81OHHMdWd6@/RX>XBVLPTHS[T0)<N,e699R(BAM@c7
J:>64D^5&Y;O\K?c1dT[bDR7YN7?G&D#(ZFI)gDKDM=<Y-9TGe_@6-GB+c,bYeBM
Be<?(-6bK:T=Cg+4#XEVFfg.ABM.f1:^d8c>b,,96TLC4VE1cXU:FWFR-JN+UC?F
WG5881g)F;0[N_S7YBJ6.#R&=8d]?f4^9@0?]1-F0?,LKWbJe/B4P,KQ1-[G:+4-
V[B)H(>Td5dSd0;Q0bf7fgLP&+c&&aDGd.VU#MC\]OM0;<;2?2<W203Q^cKNbVDY
4A(E,Y?W5_K:T+[.6-BY(g.B\4=[JDRCMNVVK3acER2(a=g2dc]8DQGVW>+?H3)V
[&.8.D58DP8RZ?0@c8I?H.<6OM-9g5PJcI4<?\,BDVDD_LaAbPZ[gSe0AbdD^\=F
aLeL=UN=Q:G\=:;J9))Eg0/C/X[ZBg&1YGZYBZ(YX46+QgNdMR,2[Rd:3E=BG=V#
0f6Jc/4>QaLXG0DGVJW(R<_d<R&AAMY<[GN>^Yc:KC);Eb-H_b7WSXbEJV9+.FI-
TEBNT@=Aede,9I&7:_K:.(CA:/9N)0^FfM^WJ7O[BZeX_?AfME0,CN:g)S+[)I1S
>9YN^#/;BG]@L8UXSASR7K0^F0)b..6cBZVF=6YEL8g2_E[QOBcd4+C=SCSILW+[
WB5QITO]W[1;d]UbN3A_fY9Q=\\&caQM9c4G>[6[PR#FKG.NK<LEaN^=5?;O&N_#
JRB5TS48_)gX#^gO0H\a:GNZeQ:?[(N1gA^ATUG,Q^CUJJSUL/]VQPQXIg(5.:U^
]56W&eC:0)Lb@M/;E&a)@)ZFT\f)8MG5/^0T&DR_eW\DdWA2PD]HP7\XLSgU/<O2
JZ\<W1Z?0.eQDaS,gf=>Z<FY=8fP,4Y^\23/OSSZ<DU_QQSHV=B@c@;Gf17=.fBJ
WE<d^1744#^8Qb;.2e+e1d1#7ZW_IR_Ldc:LJW18-d)cGeAWH=EdF;@a3b/(\2;;
V/2KK5Ub#Adb\G&5YS:Db\E0Sfd:N,MJP,)17.IR\[\3TWe]Y],G6&3cVDJ&BX)K
aI(D,<+bBHG_&:^=J-GXN81Q_C^1b8<;3S7\MK[=-U8W6b2\Gf:aLbb#ZE.Lf+EU
Dd(a0]Yg6S;0KYd+E<fPET:,J<PCM9TH0a[W;I[7]#2L45.VG3bN<RBCD]cD_K(+
P;5<<EJJg/BUf_@A^.[X;NJgNYR[EX^DR+>MI).<]W^[M#Z=E:6NZFLc2H#ADQBJ
.R?[287dH+:2GW20Bg#KB6)>)+8Z/Q49EcLM+)/7[&:_QJ8)YY(P>7P(2SQ=E\=T
V.DRJb5O]Jf?:Je7IUPU76BfU;+R@,_SM;SAID;K8;3]67B@4GJa+CEG#H1fZ791
a&PA>3^;d9,7UWe6[<<F::&5Ka.WcYfe2OeB.aeK=&CKX&=7b4K77fPT=&#B,c)6
#>KDET&@&.&9)-35/+9^HUKda>_85RbLV0B8/5FY@D09QJd.<g#?L:2U6Mf25d5g
_.7];OY0e7>Z[b42GEGAS-=4XIf2MHeQ>(gM+&ZZ+SHII._>WX)\X=.7YA\=,Jf8
=0cSFF@44]PeYXXe04)2>Y-5CG-B?=]67H[R+TI-a),LLWU3:WLS>RW?X1gGBP)K
^dTRIaZT<H_Y+@L2I&1+DJV4Z5Ia9I1T2@)&BWT,/9/G6(+cFQA27;a;9,)YYY/K
04Pgcf55T2&I4T.LJIU.[=M>7VD=fNX/,8@Hg(_+L+Z3HZ)Q?+1@9[+Y>(e)=a7]
#NBSY#E;^O-FI?X#[UbQL0Rd&OMge?\KNTO_I69b9/&H-ID.@_S&MSHNOC^fFD,N
d#&@]?e;WeH742cEYcNFd=:a^[1]=D/(gD__H3/-fOX7D6V&I@[\@R2^YF-c8ee@
W^7ceGV5&FB8323Y2TfZDV<aSf4,#LYJTL5\LNBCF[K(\AeQUSEgC?0(QK]UON0S
3,271NW9A?dNKP2&J>]4,c<e-N7:Xf[d+8TUIc27/8X^GED,#3Y0a9[fEL>LZfZZ
APIFN5F0\aC@]/2-V0O)\Vee]7[cTC#gTW&&H)U-c.gYV-VeUdKc:76N-E-Z;F[O
B#/3#?)/PbK:f99J(Q]Ve+MX.<G9.EAOF(??E4e:AA6M00(RbH5:,a<K9TZOBcfA
<8V3IOe:FPQCW3F?I8?0VcN95FYS1:VA+;IL9-,XIKLVIaJB2Pe0Q,cURJP,NZ.F
.TaBM6GcPED,]N6g^LX0Gd;eVIXL0.FRP]g5.MB/G)fcTO(,L\e4&Bg8RH3=:N1=
:BMCLSF8;/6a#RN+7CQXc(71UWRagZc[g-FdcEK^Z3D_GS\8UMZ3aM=91T-;<66J
SU&JdBAC/9-:#J;/Z>8G^H/?\3A<F73^B2U\cXRCWA<^f?b(J-:NOKR1QA@VV(TB
ZRe<N.6-6d(8Ze)W1V2gWa>-3c877CU#>5,WW>-/>[;,\^<+I6C;4/X8<51Y6SWF
F7WeeEMaK7=[OU[0\QZZKI6>Y7eT\5.VWB.33OCeg+E6DgB8=c0<R[<8L-aB:Z4+
K[),&1VQXI;>_8<43(B?eGSD\+PR?7PF+)C9b78E]68#;M>;UTCBFS+K4+e.X3VN
1MNU@JQR_(]S.5M771U3O16HaR?g6N_KGADfPE40V)4T8J)X39P/^Re?8;_?_[DD
Vf6O[RG;O]>KV#ae.OL;;U#/YCWgT29UeOU3T\;RGd8D:7=^W6)^AI8[OMW1gW]=
<,d2()VP0X)58&S[7>;^aC+K1X:+.ZQP-_61SO=1b)4-f\bXXOQ2Y4AZ+CP=R&87
<OCA0-QTZ<+9,J1X3[,aW;TZ>=\fZ:]bA-/H?JL7PZO#+MbcP^O[P3:,H.1Cc-7^
P>C>6X-S,3.]O4M-H56WF^S5gV8Ygb(c_/YS/-L^)NEUSFDV,?0T>@)E4HH1bXeA
@F@2]0GYe0^@0U;K49]^f9BbHE[(+eFJ[70A;6TL16N9[f(M&:f[TV4:#)EUK\;6
>V7E+(._<@P8HS.^g5DEL2]R.F=RPHQT2_HBaEVfHBJ\27Tb^F-0S4dAWMZZ5H<4
42C<(BS4[K[Ia^<-(\c8&d>D1Ee+><EQM;_31??VQX.0_Za:d-WCX#TMMX8Y]W/D
YC/W1&4_8[IIbJJFUNIeQ1KTKNc;?ROH6=O]f2Ze(&EE?-KY-/@64476.+;bAUJ9
AX/f=]f>bK()\+?YLQ\K>B2c/dAAgGO.YN?[Y]&MW;d2bF=K[7F7eUgJ=3=Z>bC&
,RU1TOe7N(P@E89#.<7aJI(ZdW752TI.ggeQeSeVOGOc(6?JbId\TQ>R[M<DCALA
cb2:B7D\ZYI[#8AWG4e99_[c,?eZC):IVE#B+)(;#8VV91(7F:YfADO>N=f7:gZW
KLMgFO+R;L9gMAGEH[DU=gVQVEHTR9VYM39acDN4Hb:3D[<c,F&XCRTVJ#B&Xg?6
UJ_6+JYX>W.M0<Tde^UUg:]<JER>S]&=:?K2NJUZN5F.WJR\fM#TTN&cA/#[b>A4
aT>5MN=4F@U=\;P[2Fdd7OH=NY/\[T8Y)I/X:YOMD>:KCc:#J9fDBA3(HUZRAP&J
24]&7OT1T[A2Q;Q<_I;4I+K^4UX&ed\?gcgcM1H\)G7)+<Q0FJ>)-a#OK^Rd<_J9
(?>Sd71_YE_#T<?<eU:O6Y_+Qd2>dU@V,M/CZ<,.1VWIQ4\b<B:aJ@#/RdC1+O84
85Mga2(MKQ1OMHXF/6aD6U7A\Q1gV8?>;NgVJDaYAOR9][9^b3a2Zf?DI:U6gM]T
;3I4ZLTE?U[EO[G^Ce;M5J?5aV/JQ7A4DcP;c0I;X24?>-QgGN)I#ZYV6T0(/?AX
IYVD&K/<0fS57^(d>U_D-QP>U#[1=fV>WL,KJCFMD3NI7(R1c\-ga;W3T>[1Y0A=
I;O.?0[[OQ^B>HaCA9AV<^]248:1JIe)7055cb]E+E[D\Y\]4Qeb@\bT147VO3>;
JBf;:a46;geV9dI?^VdB7-FOM\D[f(a&B:7U#>E)DTXa/?YCKIF8S599-(IXb7gc
9cF^63^-2d/Mde9\]J,Ve31e5e-1G4b/fVeBVK<KeHO4f=4I58acI)>T,&(/;WZ=
TD]XK9RAC[40U)BBWE,GI72g<F_[,1)D)>3d)&_Ng=YeJW-[P98_?R9?ZEbJ0YFg
Z@VLcO&,\Z>WU>Y33+KCe>PC&[_N\R@Q.TO\4X>_@@O2]KWR#^d?IP_9@5,I+PH<
J+QM=^,L9Pa]5N[/IU<J5E3ScV^V/RQ5C&(#9JN@(^5D\8=AUMb]M[^NfGdWTKge
KY5#a0_N^&c]ARA5=(AB3ATS[F4P?c(^Z6_;3He8<b:=#]K5G:Q?E.Oaa4I--eME
H(\H8:\FgFe#89?gG:U5PcUYVG-O0U8(,?dNN9daF=;)/<:/fd>\-LfZ6C2XU6Cd
<a7Q)<fZ?Yb+S;-U)<T8;cIc,E.4/K^4X[)g-9?PD)7&K7EJW8KcVf4T-3?TB6>a
A/W?Y5@<B1B=;YO32cga/HW7&\,KDLJb?-7,)d@@3<,#(Q2Q2<LcPCGAReZeXK3(
3g<S(XXf.\bFKH_9(S_>,HLNNQ69ZU@0U,DP<_(dcAH9:\?eRTfNab9H#[81cFAM
\CJ;b=07f5JJ[_64RA+70#:<5(-KFa6A\#ASJJ\@EGa2UM]973B@-5_^=bc4)D:6
R>41(TKc#1Y3L1)1#<\YR,#T_N?6?-fOL@e2-QbP\<R)ANUW7d#?Ha5-V9,MLH_H
951GRJ<30;bBA.^6NUa\#[WB7UL&@>QXFa=_)fI6/NBT,d119H]5-CAJ/g::7dT.
&L,dOU;(7(.KS&\JLFMXN#OI4]ND>A4UG:A.,g)_3?,W-AW[UD7J^RfbVd?)MYVR
(J(_A93?b\7\bbZ.?)KW\9421KUT(@=50FE9a9K+Z&3.8NDdV:Y3?B_.-3TJ16RZ
b_498.\B(YPESeg^MN71+DIe?2>&B\f6.#Z&T\ZcJ_]dDN)I-dQ7adB4-J>2)BE/
XJ<POY_08bW<;4)a;3eSK(6^Y^Ia1Z,?=d)99L/)8?X6@XK;-BYf9+)C4PMZ)/BK
3ME.Lce)<EA9GG4]8O_CY,>K&O@=d);P&B7)WV^71YE+^#9KUWPf@1=BG4MY(V#(
O=SPA?P80dBYg<B.cVENV9@\+g=+2a;/-&_aXWfG=>dVe4_J6,fPWFbP9\GeUVRJ
GLVfA-bJEFKAcH;;J99#5HFR1G=Za7GF[Q7YN&M+303(__](C]ETU?9<52g8R/g/
X>FQ18K>&d[Rc&-:@Gf[2S8,/;aT7-M&OB<eO?<eV[1?_5Jg)N;R93SfcU9]#)7Y
caAOf&]L,8.?XN\[JN>eS/[8SF3)</#GN;SX-Z<JZW4[WM]>I3SEG\G/X+DEe\&L
R>UR:Z+5IcQR\Kd0G.DA9)06?4JX8CYFJKcNJ;-YHS-:g-\a?+.c/:\W54NK91dH
KRB@f/18Gb2M]7?HI9Z^A:]4FO0.G5e1KGI>_.^eJ6<-TWZ._2bQNNO&#?>a;c07
THdF1a1g>-C>RI<AJDM=UWZdAT3/VX2gU>c.UeDN?\L3R6?a/ED[MF,=dA;0:4AO
#@+2&.cN21[E+7?MgEFYI.d,N0?C=_EQSNbRG&W6]05Q.D.F@d.=;>&H&d<SR3HX
NN[\J)?\Wf->8;@_Vf\SRc;.6NdBfD?XgfQbKRBHNc/g(cSZK6^S/GNa1<(E4Gbd
2bG4#94&4WJGYYd.YFeZd91<U1SRL,(F37&)ACUfM>3ZOV[@d>GZ]OcC.>>^G=FT
=M6S4]KH23>gB)0X.:UWK<+W(U&TaJB-<:g4LN5f5EVH<T4PG6bd3S-YVa:JF4fF
3(#SVZV[VUL6?I&B>3&OB8JA3G\ZJfQ.W>8/@B?XZW&32:eCeK@AGS?\>37N#E77
K:D\bg?:^PY)I:JZ.IXa[4b106CIQL8N.:aP6\;GKWA[-B,8ROS-[N,/N;,1Fb]D
bN22Hd9ROA),egD@8ICN_>0MM/\^Q<da,H/W<dEF:FTUbf#C=,XPI#K?d(4b=4EZ
3Rd_E3?.;OLW5HPDZ8PZN@fCS-1\A<>XBY9TfPPU^M;>BN1&RA+G)6\G3D5/;)16
e8M#RSQNS?9;#CF8#).6CN+N3E0L2)Z79-=F7<G(D;#@#?](FA+?[b4)]a<2[F9E
d.R[f&FBK(b(EDSY?3Z[MUX9(b=b>#R8)55VZ<CUVK^C\Zg&a&5VTXdW0?DG&Z#F
Jf&[]QG]@8X8J?9B0+,N?0M55;O\U7.T>\aR2Q01ac1DLB5=8ePBN?7.V(fV12F1
K48WCcQdN6&Yb0NZYY19,P/;#AQL\AN#GZU&B-/,YJ^V3O=,-ge.8Sd@-Fd1R.7K
ec.YU)/@N@g5[;Icg],7TCEDGGAUMSF+,/6Y_&,_2#.0VBV:QE&KMO#2(<82C5fJ
I5]:U[:MP6>ed^c[NP>G5).LQJB=_Sa_8B1WB@_A>@9UU^Ua/de_NNGRR>U-MQ\e
<^-9[7CHSKV<\[YMSd1P<5LMZL5&9R+/DS-ggc;a4)?MCM1CY8\6D2][@WPJ)G<9
0)\V021Lc-7V/#]1N97=/Ga-=@[.XZ?PM_3E5UDTIe.N&QJgFP+P)RW0TDA)C]C&
+<[CY^PETId6?/F:)W\W/d_Z\F5Z1T_[dK]QQfN<X3UL?YT,IE]H_&dDA(JI7=P9
QPG2XLN]fSY\,E,&fNJ[.J07353@4[)NQ&J@[d2KF2U;35Q3VDU3DKeP)8cG6-;]
AD>ID,6g,W,D+<.P0E-\,:Z?DU<TVX1A[VLF6+gOg1U7BeIg+NaGGZf>(-eD)],.
\?fE-6V8e86R5Z&;]S>EW[Z;69d_&Y(,5-0bD?:?010:#=;(\0\Ed_QE7#35OB<0
4?(YG/E,]&(2,cI-S@e6J8+F#cV+@<ZE1g>/(0YJ5&EJQc,NFX&LH=9CWX;f?[G.
1)9/BTRP9C[KS</A>&I8M0V2PQH?4TPJ(/[d(D_F8RD^N20^?Od\.VJY:-;/=OB-
Z9E&bg#Y=c,+<Zc;LH?8YGF6R;(QFP<19#>0QU)^=UX8]NfdQ,A6EcaY66K<QfDc
&9Ve3B0EKd,W3)R_1;&:J/0IE[cZD=A^a>NTXP>6]1[/+e8(&VZ(7D40LH2B-eI9
e5FOL[B(bK<8_E82:2PU[Md;aTY8\::-,+_]+1)HL))A=1c&:f?..Y8cWBP+-4gK
I79??5;H,aTHTbQ=RFJ+f^_5Y;>\.2SS^.DB52[Z++-@a^B0H?.JLNPf\MB^Y&CI
V/=[YYJKUGX6YgVgb4T9#Q#eLT<WP-@YS2<d9,f^_;YO&W-T3;>2V591:0fcX5R0
+??Z^\\.dZD&e8<WR[@fdegR[ST5C-)\=0a>H^WIKZ@RO?DN?fB^A2\C5KLZ3#(J
WB)+O\:?SO62\].B_B#Z?bY:+)[7CCH8Y2I5Z_^X\^(eCgcV:_b5V<PC_Tb2ATCg
BVRIb#)4T=H^3I664EMLRc6f:=WeaR_6^FY,Z80)]Sc)Y+gCU3@[Ed_5(<AY/2S9
U8^aad6PbJ>0=[d.0M2PYa=[(<&[b#H[<.B]+OYeWWP6b1La?cN>#+f64c3@<gUU
TCHBR/E2@6_4YB[G[@8\8#fbH_KLV8aM.\^18/S-\6QbQJ1^\_I>@:QU)O2RC](-
LN)AZ/;+-[/U_^LgaZ,dA417)>Z,a_g&/[.4FEd&S/;R\P;5g6e3]Tb=(TEY;/VA
HFbDg00PG:Le72L7U0#8Q;:a&Y[U^S[:?_7;ONc17&8-ga,F6geHcB_+0_<,\@R_
g5a?7+>)V[J/MY(70V[4_QRGf>.V418Vb&4=VUS0H.8MH,f4(Y/gXN:=f;1H6\&b
=f.P(R514OD@^Ge+dDO\9R-22_Cb.ZBM/D\&JedEL^DHOe3a;[=RV[?/-A&WSVF=
0f.#O=25:NJ:.A,IW3;GA?5RHTY.6RI-7H^(,.OO^AV@Z)BaC]R+3g1W:?<\&VNg
;#:fALL3]2388W>A2-Dd#>--@FCEQ=g]2;P264,MVOeHERD]R?aX\=/32LFTb/\0
D_M#f7\]C#g9&>@CRHdLNf<&+Y<)ECQ-d/L:g_e@O?b?<?3gQgbb]^AKHQYH1K4Z
#_7_5D;B>J1WBY[]KJM+/;.DDB2N4PQ/\-.Z[#.G<3gRM8<2RB?^UC4D/[bEB&2?
.P^KbY^MX.K34S)YbFO4@O6c1?N6T)c]D_/\<Sd_5YDV=XGBg\,5f9,A7(]JM(F:
de/2:.DI_2],UJ0VW7X8ZY(2G6gEdPfB8C;MTU<>]<N@V0]R/W:>;JSTP+K4La9F
65@eY0?dJB,GMgO7DFc,K;dT^;CCZJL/^=1TdHL0R@0=7-aCKJZf_)TV@:TS]QK:
_1/cLER1#_J;aaCe(V0INf[a#fF8[O()W0_5^R8gbP/T\;2A+0T]d39@MNdA2aBT
3(ZdXa+/QZ@K_SUK/<2H4LEQONF;2R:Z2S/X;WUO:0VOTf;->-/71?Vd=gHARfVR
DQE;.-@CbMWUE9fU4(BVJ_=+NbeF9VbR(=[IF2@=CXV3RNIdC]NFA5)ZbgOK-S[_
40PG_=g8]<FfM,M>dG/fGEgYT?]X<ef@W48ED1J;7(26IOGfMId80L2E(F]MCWVM
Id2X&&#U82eE(76d=68)3K<AN]F>Ea+bIC)(^PI,AZM:8)L>/c+).(C[1?:Jd:6B
VOa)]3R1NIOZK7&>?ZI<3?D2ID3DU42g+X2[@4ICYXf;)[F8&7L,8>LcRBTYf51U
7<?HE,@W^b+&a)=C):f0/J\BC_9I5?^.LW-8+H>U8\1@)74P<fYE-1Ne^@]-W5aY
]6-+AQ5aM[;dLR??O3RU/#^AK9-D^6QRR=66KK/=V3O\,.(ed42BS<Y[=g^ZgfVW
FU9&&2D?Q#<eN0W4FCHH.+JNCTS.c_5&E)BcGEB6@)g]Bg-TRTJgOD6XbC:Xd5[e
)F0Y(5^MRIE_(eU+VZIURDP6D0XWY&Vc,&GL/CJV&U1M\+\BgdT^baDHH>KUWf?#
>HW[FK^Z@IWN\()](Z838g159K(7dUfdNVJS>Ega6Y2L7IC66>NDOdG]BW_cKJMQ
IBc.DQW;PLIW]N0#4Nd;-231+9^4NJg+ET81(Nb@b:M0#E_;6cP1ZG:NJ98.>e)(
7b+LQC,1[gW:O_,BA,0L_.IT+401EVY3#DAHGBa]9K=Q+?F3K4XdD:RV/FC_A1.E
?ab==O\_bQ4?aAP0,8dZ,.,;?U+>.)C>51WZbD+NZ)Ca[(G0QU71g&XVb-J#1Pd8
4g+O(@S73e@49\c,1B[.N@L=,PAWC/AHSN:MRU&@CcdUD>R5,GP,8;-^\JVbW9=_
05ffY>+/R,[9OR=68U\;0Z:OLJ(7WfP)6X@\cT@E<1dee;^,UDEPcCcGZZEcVC=&
LWOWfRPG)/>a)5f-f8))dWZC2R=BHM2Q_A7JYJY13-e7@FXO51NIBMC=4fZG3RdB
E#KB&R9N,0L]2X(DYf(7cYNKW:0@_ZaX<B=fP#b)[\FARCDFZ6c]WQ>ER[IDA^OS
=(5;c>Nc;PCR&F8T3a@VL\_=KGI?6=Nd0OEY:SX2]I7GL^5[ZSXI./:?>1?/<.U]
KA&]+K+@ScADCI0QKeX:M4S.a?gL=cbDf)2A_7O]2]\?\S[[M-?#8bS(XFO4dOME
OC<gU7GSH2,g#@]DCe)2Nae@>>;]CG-0K(Cg)RScTg.0/>bIRVd]0D\;+Ab+c5Z7
8dA^#V4V[9-N>ZNP\6)1=YRJ(UTS[Od)0G>dYRA<-\_.H7G3aRWMWGIK<U1ODN2f
a-47\(0X:+RE&.>=#HQUeaR(2SF5HL/=C(E]EJf#_S7eJ0+/BPEW3IE4ZJH,G@Ta
BG@;Y#[X1_:_8cH+]^V&VL>gOW_I]d49G@VIHUG;CUFZK;8e:U7-;3A1?F6eJ?C>
44WW.W)5a-)=VP&H_CBBRe6I5V7H66=ed2U-S,f>fG-dV>):H^(D)IB@WC3>Y@:G
G7dGY=-E3QW(EEZ(9N(9+XF0C<)80^)=:cbM0SU[=I0B@aZG9RN\<b/F):\FW:T?
86F/Vb1)]WJ<g,:&CdcafJa_Mf#^PAf(S]^D>X]9(fDP?TN56Gc.aQ1e#XSfLG/6
aOFfa))aX@C=+5aI[;@OMCL;ge,Q2<S7\bge66aGWcD<J0g:TO98H8@:CEHZ;a7/
H(,fO\K>JZWT,++Ha\_b>Cc2bgFC>G?Wa?SD2051/#J9F1MC,A39f@=cc0J@)NZR
3ETTLVDZ)9+;O10DL]edXN^bF)+e:Da&YYL:3H8I/B8WICXMN]RNO7#b#0I/YIWW
1A)5Y.UC;U>Bf#>O<UL0CZ/^4IY^NUa+2g:?(.0ZUH3O4TLRS_6c^-BDEF=5KA,d
2&Kg\FD26;;f459:Q61+_d<4LA4+YHC/[#PWCKg2J#AM[FSNW]]bbGEaZWM&/7f.
B&c16-\=9Y44YgK?J7EQO_/b4?GP_OG-H5T^L7JU/(&?(AVTFU7V_b;>I5D<F(9Q
3a(/_GK-S[:RFP,GOd.\TN>9#EK9D;EY/FRRdQ/J?.4>Sf[V7aMc)8bV3W1:O6F&
a;X<+2W^XX8KY)4P9GH95@([W]M.V/.+LK3Q]e7\Y]aY;Q3F9-HJI^>S6->(3;F&
M9UZ51\)H2.?2W&-R^?0&eQDb>/Z891e<^>\2KU3b=SJWb#V^VSIEL7_/BP2e=cF
Q)=D&Zd8UC#=L6XI?EOZ1\Q2G?V<G;b/IP:^Lc@ZNQ(O?P@9cAI,gFfa38WR:A\Y
YEaBHF.594018:UO+89M>-@,QQ=(<Q5]HRPV+ZF/I>;+QE#@E9HVec3BJA9S1RE@
c8TCN&_P[KFH5B#Y:I.=MWHWB<24=6/>[R,Yf71).=,Hd<Y8B9V?C;+4FbIMU/Cc
R4RaT17AG;JZ>6,=JCZAQ;LEZ2.DV?NB@8IC,B\G-LgAfP4MF.geQBa1EZQEUR4P
X&/-]PcXN^&+3b>I+G\9<G2U]2gL4+ce=aQU/1Z_H#M50\A\8eUT-2<=M\Q=LZC]
(+BH/cLKPS?Oc9Q@FW@Vd^)/KbEf)KfH),SM_I;d_Zf;OTa6>N@?WGC\-IEBS1_M
8_7S7,/Sd(20@QcC.IJ0QW,dfXUXJ+cY@I#UU_]1R-+YOe,:Ag=[^FWCV>b&NF27
)@?JZW8?=557)N@FC<_U[=G@NM&Z34B_;c3YL-dZL0?\D,>\YC^#g2.Ce.0FG<6U
H-W6)3);6JQ/dN;W2]W>cPZ8J0^JR?A9=e[O-5SF6HD0TC(Ec]?-bT(LRE/^<3MT
99F>IDC#S(C/;P#/a]PH=@W66g>)]e@I,JL#bU5G<^;6YPZM#fLdB2_D8M]@]_C;
[:8C>_H6H1.L&;C-,&-_5fHfZce-^#@P5Pc&EV=-DRHPUZW5Jgc?:O#I>SS\&ER_
ZF3:Fg&/Kge3\g.FU1^dcQOKDg:NIJ2K:)Z>301Je+],OcDXTf4XBbZcCS90B=?&
6@He.3;3fTKdaFBLS-fMX_d5]2C)W^FE3897gN^#E_0ZZcQ=ae/8C#^8&Lg>^._Q
L=?]YTK(FC.@8]_8L13/MdM;.Q<1Dc?5<;g0CL;aHB>V6+#KO#]X[R0<Z#MfR6Kf
H54EX4GDP&PRX;ZMH:U1+3JYWN:R7F&SJ)+]]^[GQ295@EO,OfZU6\Qg5(#gUYeD
]Q]5[+g?;eB+O,[E?,:QP2@A7\59X]<WXAI1ZaNKORgWU9<SIbFBK,DOZF:WIP_&
W0a6N/(f2@:Z]NYW/OYJ:E45.C-KQ)7>HI>b^0#D;2HT=9_>A1E?6MH@L[;dBEWI
]R3Fe5EO/G&5G0=9[C2\G:^7O<HO2OM.PW)1-TU0.:MOHYH^GS.N[;MVfP=04QDF
#JVW.C1I.+=I@6##\2]4_.E-<6:Oa@D:]7MeA[ZM&?+Wc.S4M9AG/Q0Ud2b<^eI2
aR,;ZLd2OIPF10@g^VSB1+>)3JbK??E#b<H0Q3CAg@MbH^;1U]]C^RXCQ@<A+TYH
/O=3F.B<Y0G_<+]JDLDd6MGO&1N2]LYZC[T\[g3JfPW@8STg6>9V<)>UKDTHE<\=
5>/1J/&L<?c??ec<(D?M>QE4C-J_cagP08&X[DD(^QPU>/6gf-+CMHP=UZ5EU/b1
X8&.+>6.DIG&7gb,X[RDB7OH6YQX,^M&\AHW\aKbY())UB.Z6-[YU0114[?@=LCC
a(&b@:g-5M8_Ad39KI+32G\A:)LVJ+O_Y]Sc14&N?09U/,/57E.MgIfJP>ANgMK=
4H_dS-4782>M/<F@BA6(,593B8=7)YR0Z)eHHN+g2P/>@\G,(;Z1#bA^J3=e(NW<
N+?f2\:c,GKf\2^8[:#a)-WeJ5b0UB99.Je<;X_G[4bT;ggI.783/b_G,b-39G@^
>2M[)GV9L,9P^:AZ7G@V;Hc5>97T.?&#SOXSbUa--b6<SXTaR0ZSeJU]J<2#=CX=
DO+\QEY)Ce<R?IP?2;SXKf@++eGJD=6GAD91.[1M3V2IT[?<Z\OddUc.:76=..dN
W7cI0S->fW\PF_d/@4FL[]V38Q)#bI0SW-[NCM5WIP9[Ze/9/AJ;;#M,59e<6<C?
X9M7(60JWD:,/^(::FD&\4/,8QER/cQD/@B8M]=;bfIFV[L(,RB?2P8JG]+gY0,V
Y2;))-IRUb2:RHG/?&)HdT9\1\N3RLA[O<SC>f6,>EcV,9GG]YSZ7;XJU@;VQ];b
0BT>M/SE:B+Y2>]<.HQ\d,(-^>N1^ga??&J):R;G#PP:4==A\a5;,S\V+,:<3SH9
\\S\d)YTef1[FMa=@bQ8PUAJ4W/C@@FWFXFGOY)_+GT,2YLA17CWN,6)UcKCcCOI
GNAc-P9F=6E&;9H@>,0ZIP;4QW&&AK;8Mb6D7g\YT<>Uf^Mb=/gZ?0NN7>4_\aV?
RW]DB?5XeBHB8T]S#K^?H@fXDg_3R<-OFe3(HZXIKa,:5fa_?6N63&+PT(SgXWOS
DV>g[gY<P=gN-?Sa-Y+I:Y#BP.S=?K&C+)XOOB-[c^>4;17?>\ZdY.)W9c[2@e.:
>3B/Sb7\f\2C[S_8J>PNX2FL,:Y=XND6g<4SB2EW2MfW[>I5\ZW<NNW55_QW=-H5
7R_(B03;J0XVZOeR1e.XW+95b^)9:9ANOWOMQIb+IRA&R#QIa)=QW-7SS;6L;S:<
/VT<-8F6DU?dJ7<M#Dd8UJ^PG7GUJ0a5YB=?PNG]VPWG[KFXXM^cVER,JY>6/aXd
MS8RRM)1OSE8dJZfR\86b\,WAT9&g)MSc^8B2^_AU(KA0daR#I-0XZ?-.#c4eG70
KA<511VM(PRH;&fBIK7V3NQ_W>g1#7W,Igd<+2\XD9[(8\#3/1+4FaW5K/8=WEGR
YA<?Fe.;=R[68Qf8E4b0Me([KC03gg.SK88b#+PVKCU1EVI2].;.+<2Y((:9^N\(
5g@44+F\Xd11ag9XQWQU<Q7c5N49]Pf9A<F0CQ=7=WdXI?--2O?cY-2H-ZF-c5R0
]?]+4W3LgS=HH+\3((^(K8P)2L90b5T^.bKM)g0T_T(K1=d>[UT)DDa+Z4]N;Yga
a>gEae7BURJ:9H.QBT,XI:S_eJ)NbAPbYTB&cR/[:J0GS>;D>5CM@WMJ<:@&6UI]
2PfA\K813E-RH]FLaJ]>?edRKH@P@+9-gO8?_Z[Y:VE/<VN\dc(_aZ4SU#KNfR-R
fQT,&SYKXd1/IJ(]U-X:+Ab)@7==fLQJA#dK-O^0?W]@:>5Y&>6<8f+K]c/K,91@
VOg9MXJGO9+\M/^2S3E#JcT57^,:7]b90Xc2[96&7CUP<bGXZe\5?VIfgZ0T4I7V
-I5))-e(]+F;0e[(:J-UNC0]QcVfQ+&-eL5/A0QT^B?Uf2GWCPI9@TNL;Y+9Z8W<
65eX1:5M[G(8^P6-2T@<QTf+&-/e.U_\DYDM8)?^/OT^8/16\R;YYQ(Tg_E>J&46
aY_3/QF2/)Q8/+&=dNN6gcWPUdRRB@(f(2R/H6DLMMQcQV7N?;ZfOfabS6GFU61c
2d8:@H-F&NF9Od#VHFAd2;b4)WA2=Z1@F7C4DY/V?02JG;;e#e)W;+S&Y0_[9EN)
P\7?g0SM;P+C40EY_N5:GX1BWc#aTTHCXJe<fYUF4.-FaIS0QU^&8@c_N1?0dTIZ
(Ef/0P(WR@&3/c:ZBPZU8_.:\>GP0#:L0-B,@cEOQc9S5c93D^dNcNa.:\>9b.?4
#bcC7dSOAc<dST7:[P3QJ;F:3J<(fFMf,?2#1Ud5V\SUdY6.ANbXYID)=9K9^TAN
PEfZ59?;YFRcCeXb;+36IK#RUEQf?\-FO:_Hb3)A0[XC2H5<#b1>E]?Y3c[gcRW6
;IW<GO2^=B-6-Rf@fMH7<33d#Q+3(<=^/[cJ51[DA#a7>4761V;]W(@(<Ja4)V8f
MfW6-Jc(:R-^,X7,[e:WEa#_eFOgYLOLDL<(Td#SG)^)^OA3HWI]4BK^f.8?KQ=A
RHN?+C2Q]Kg(@7N3+;)+5:P_+@+W]:B]f)dN9E1JMPgB\I7>J;9^>\D3,6S-VOKf
[:)XI),8Q2B/GGJEe+X0[7I8W,b=PcB_[62N72+4FQ9YEec#J7L03gKEe:Xb_9[b
b[YNYAAK0f^G(08375Y,_JAC-Td_L?FO?E.FLO[Z9b]+\Ra&#F9?PV>G7<LDf,#,
N-N^gHD0,K&448_&OUW[-<Ng[Q,e6_/NC=N/6FaYeeQ#,H@WPKKaaD<:\\ge]A-Z
c(Q(Nc]6MXd]HbGSV#[=4b8SS-V-6]ZT=L3?:f3@g=T2:Y>\<^He<(\C@^D-S4)V
R6F[TTCf9^?63;?&I0=KBSS7c=c@0Q??_fNYdM489Tc57+G_)>-3c-RfV)WC-OUU
KS:I,WG3)CX+QR7]@bgLb=ZP?PR+IO)<eZ33_L]F)ULSYEEIe:U,57OI^C?Q\Z>A
<7,aa;_0L&BgNU/]-3Tb&S/FGUQQ5P@BF9C?H.;J)4bc&7H^R(-4Vf76:VSNNeZ.
-:a^2/c@QKJGI/4WZg:#R/V8fb79N3PHEbC:a1[G-8b/0>Va]0_fJ)=H-[D9QS[b
gd/MfD6/3^aM69F<7DS]a<]X.O[^GU\@4V7U)_3ED+@WSI<6baU(L^:f=I,0\MP+
(MT/44)([@A26F1>KS3aA)280g+aT/Q-a&08DJ04;:BFQ6dT^[-;>5G95=EV2ZJ8
cN_HZ/aZV?A)NX6?J7Ua1b,UM=[Kd#5>bH;>+G1W<b<1A)8K^fOFVXL+DF/A[C(Q
J[E>(@O=>P>a[AY>AeaQ0A4b6fI(1D^2;Rcd4?\0<,+V^&c3)A@J^SZc]-<GdSR_
dccI>a2:XLDLWgMZL\@5dXC1We19.#=2E&G:)cSf1E7AfdX.W1,gRg/3N2ZS7eCY
;1)=f_\<\JQFCHY?2PGfc=>f0S/I]\PbefTW1eNJGY0eQ_D6.7\c.LKO2MdFU\\1
T8]<FCa+VZ80FN(+GX\_<8G;6I(R5NS?)ER?Xc)8\PU&+_)HB:E/4V/+D]MA;SIJ
_fS8O>6b^N]R9;e23#^GDf&5<LSFf/T4,OZB<d75AKV9(QU_c<bWNbc=bLLaRZNU
B,P-aSB-3;6KII<7U4F^b]DXKXXCZM@0HY(0TSI_Z;&Y=@D_^Y+dZ],Bc7?YGFOS
.[I3WA&g)eSW:7cOg3F@..U:M,L,>bM809Q+::A-&9T6H8bgg9T]O^Q:5E,B9_9X
g?787TeT\#UYPD;__Ag+;7RUM6+SK#MB=L:8A=)RRIKSTJ_;O8I.7_M5=^=:&>)9
KB7PMX9Z0g+D:>:AU?OY1,0TK>d0@I.KK9/F6.T^b(1UW1RT^eJAP:N6#.T@b]Ge
)RWRGI1Q[L8ORR0aB@C]9<:IPGbMH4gWT3+?O<cN&>T/K,-a4Tcf0^,?-1@:gPTL
S),<d)2IOA_LS7.cc7U3(O&W_&Ee?6\27Y\;TOS.Sb]dS0,RB>+-JP_R2N]HDHF/
OQ<A,K7ZB-SYOe5Cb)2bMW;<#^X)N_bZS?Y3F)[+E4=_1A.8_.J+eD(gAMY95NT/
TDAf[B0>#WIffS7V5V-H^0V#)F2bG_N=Ob:S0DKSKY::H#_L2I/;I7/\8Fa&NXBX
J/3#3BDAgY(]?P,gREG\EJ4G4T+HQ[S;2c3J-P+.3^ER#@)_BT4A-c3077baA1+A
+gO\\<d#FM1U3:Fc]52;6MOW6KO]I-:^#M++^<TIUJ93KN[ME9#+Z_F&7[:d-JI:
\)XV+7E5+d?eU?g62)fJAbJ]^1fWc-76RUI(_^8a8)^45R2d[_C.2<5,J5W,aMMc
U>BBd^MbfS;GAZERVNaAbN0YD&6@8BRPZf<#&-Wb#U5E?<)aLOME^YQD+6=)EV[g
Oa25d@De4^8@1H8P_=f4JJ>TC;DJF///&g^DeGNC\,5MdR84T2<?7]LQA0=22JE2
7e]a8=C#9X.e?CSSL_,/HfLfMXY6J\eMLFEYT^:(-dSaT@^dX@,>aU<;P5FfU8^F
;.N0a=.)0;G.c[8>d;;]XTgB834Z;IUSeU_c6/4=#6]-^cA]3\b)c42<P3Cg7>M#
Z</O[>IO-HaJbV9Z[B:9G.TY7O.\,QF.44B^.3GbgKbV#NUNLO6#L;b:E.ARdf&-
?]NfG4XUef9gVRFT:6;89J?f@,ecF?FbR3Z9^?W5\+aPZF;.FGe7Be^fT:9@dNdJ
+B7(VDe;5]<JWKA-0Kf1W[:b74bHgN-NeaK#G;+L8+g(fS+(6g\YgVB70G@X2LM>
M0>01f&If-=ba_09?7/Q3dA#F58<d1g@^YN8E&G(c4<IM#LE^_GU-&#,c-8X:Y:0
WU]08dfX4KI<8J+)@I@84;_0/8bHHZDJK)(RILYS;V_(J_ee9CgP_U.4&Q5.H==T
/LR\WXR:b8+Z2-#LFWWOVc(E2@AXYTP8G1Z&7=P\e4L=,(H/Y?V/Y4]]Ld11Y2\X
d[KN(LPLfP>>4?)C2/=e_cT?.ZXLc;fFSU38.K_H^;8e)]KBSV/D@fH8[gWQ_1.]
[__KXQXfI@/VYCEV9&bMO?#aLN_E.?MGe?US.3T#MY]VGLK5<)0?3JG4A7_MA\=^
0D+f/KZ[O;D(D@cM9/IYJAG[>W3U(LPVUE[E[T(WJLSFN&)QOO^?AT6B;(?g0d+X
M20.Wf@4G(3.:K+..Pf&,dJV)+M03-Wde7KUIBK>J:2#bK6&7Vb:SF]SN2.6:b].
KXPTc^+>23._gR7YN\+72D+)P<6_CbWN4>:TZT^J#YS5cKLKUB1MMD4<-KVe1K0V
Ff4Z0PV@HC,SSd9\GeO;aH2-?4Y]/RY0G;&2:V6)I2?792DMUNd8E;5c4e<7_CK)
>[;4fJd6</-UU\aPX?()6FN<[EF)I:]S7B2474@:[-@2_5b>;/DH>XE>R7\<.2)/
E:;UP@)OX1G\SbE[\JI2bY1SIdVg8DV&>a+N19gD&+1]M1dNV8TR.<^<gd/[Ke]O
)O;c;;#;\bJ)RbQ^^Ae?UW6&\10.\)3AJ;&G=f8SEAE&d18eQ2/&GFQ7JT9;c,9F
6Je\H20JYgPLM5L(K]4VMD75XO+G9/PgP[Kb@_M(MLb6VOM>B;@)@[3>C91FDA+D
V1YbO3;Y34A9FJBd>\<V(HQb\,\aIWcDUa6CI3-A@VT0NZTM?9]BY_80@2^3ROR#
N_9)]EQge7bV7Y,CR>e.Y>c0e..8QGGBT&Za=?K>?6BK;&=g;f=aIgdKGGg&RJVX
&<6:_9:ALN596HM^LPL]BH8MfDOQ\5DQDK0,851?I\EH3@WY6_cSK;:J8:PJZ#8a
>RfE_+aAa/,G)V2\YE?;(2g95>D5O8.JMCdS-F=_KF,PR+COgZP+DPK8c>?U:2JR
8:KA>b<?eZ=999[A<.ObMf&ZT-XV8bK+0?6&5YgC#<-aYEc-Bf/FJ>DcbU(T>GE)
^\)R9/@V/aB=G]H)DJ:,8=d1=abFC0A+E&<1D=Hg\VG_\QbfKHJdLg@a9ZV7c.[d
#F07e[eT[+;6d#6\gV;B+>Z(V,I6Z]aV849TDKL7e//XCc?.2?3Y++TSNQK=2/+4
L[HX\I^2,[F[[A5<&>[B8^,KIFbC2><c#>D.(a<FOHZ55R3/[_ZV6=8Z3;J^/^)/
R?_9U8P7S<I,MU[1A]7#MfMY5O:be\5LDCZaWPCeM_DIU1XGZ]^a\?+]V[^CdNT4
D#-]T@9[;6,T20M@dC>;6]Zge=-cK\7F4f<D^=#?FV+bBRa-6@S7R.HUO?:Y3(Ag
.Ue-76:G#I3Bb14A]PbBUNK:4BRO2WI_3L[[<6W^5_?e<?)^:V+T73/R.M><D10d
9R68Ne4C].Sb@_5I)dE\LD]1PO9;2_FIYY/=4c(2T=E)4GeB(06JEJS:ILGK3Zd6
O3-U@0>HZ],T6YD-LSg:4S9]H]:1JF,_/T6gT-H:YXPVY^cN5GbN7H5c>]F6J]RP
.\gPSCS[=7JAQa&c<-I5d-1c\cT80PB<2W:AAUK7KWM(.VZ^2:e_,DWTMW<)Bg\^
2<d56@J:;gZ>6=[@c]W@cR>?;gC(.P:<+<6PH8DegI03]=00[MU<C]UW(1&N#Xe_
+B>S1bH1^fRR/2,@aaHU:0WLT?R&-VHA(2+F7AM\X.GO7:/_M;2[BFHM3-((]9Pe
D=@P58>B8]02(-EFda?5KeTGGT,X^GQ+;]@<_E@AJHX-(?EDJd?,V&V#F2=^BY>:
M1Z&SO-f7L1^W<DW@XK4Q]Pa6?R/?3V<[9.8I1dAZaV?QZ).@&8U9gEENfNZ^JCP
(V,ZeaY^3(a1eKH,A.e?Z0:<G#ef?;(e_0\DgI\I^[Hc@K>2[W2).L:R[RT=c=6H
CZHYAaU?XPDc&g1aMN7N@OI_,J([Hd4&<61[FH7&BW/IM@S82(a84<S]2VJDSP>G
/W+,<#,/-g-?UE6K3/KEOY<JgcgSKI6@+@0IEcW_,,S8;=fd9@//+=YSP+30H=;1
cW9,<YHa)C2KOc._0_\2P+_+<@<0[Y)DJW2VEII#.2V]c]FSH=\H/J/+-#?TV(@S
aXg7I-N;\[gN6D>&98QP@>)TcJ>BeFcI_>cQe7^U(1_,B:-7#[,Yc)TN[)f3.acf
GJR=SYV[)4T<5gJMf8(<>.CPE5:CP1X:ZCBCZd((cOCWI06=KB?_BU.+OgIc+Ld_
9=VF2QF?McARBb6M8B:UX<&5LXJ\@23Q?)G(9)d7.N251@:4QL2Ya0e;T3H.;E>e
Ld-@_5B\J,W^B<NW1-CH&(/>f0P0H=a1OV>2\1TQ@LN74)XeV,TGbHPK<2.Te8K>
S[;He,RIbYCV9\IGSf:>K7+4[D;?<X@2Z[CA9\Ve7@:Dcb3?RPS#(DgH=&&?f([N
IYC+e,b&(V;(OUg7)49YJ^T1^7?0M,Q>_dL?B:@aKZOCVNEZBFQH>1L=N+FIFV3^
fVNGTC6XJ.gILIBD;(<EX9#PFO[2WKGb+e(A3\.9NI6&d#PZ)RP/FF\LA>8&QY9_
[RB@Q[J_RT@C26HODJ0(MT^=[/aa)cfaO#MfRIZ4bc:6>_E3T6eGR(&?8MFa3Z3A
9)K^X9]e.#4?N>G8dJ:FP0TX+A7RXP#B34MWC;PRZ^/K:[a37O+^20MeAQ_#\7\=
XLf3F(>,Fb@f/d/,;;Y,1TWKEDe@H.[^a<@JK6(9ULMJ7/S2I^FaJ<:RH;+H0@S\
1\;XP46D\eJ+3=S#K:9\4beE.cU9-=9dQ&?AQKT6QQ\E07<7)7;35=+.egJ8B#P-
3Ud@,34]F]S\@#3MgM&G)&.73N]HL]7UAC-VVT/9#[1P#R_[7>L6D08(J;]T#B\]
QVX1@DTbZaPJ+a/D-;L1I3PCa;LE;KcA0MgQ_@N:ZF;70]J)O&S=UG]MA@M0GRSg
(Q:Ce@)WV6L\]PGMELGB>5Qde,&J(6<K:e.D,SD#HZ+@a?fO9]C&53]ML$
`endprotected
endmodule
// for spec check
// $display("                    SPEC-4 FAIL                   ");
// $display("                    SPEC-5 FAIL                   ");
// $display("                    SPEC-6 FAIL                   ");
// $display("                    SPEC-7 FAIL                   ");
// $display("                    SPEC-8 FAIL                   ");
// for successful design
// $display("                  Congratulations!               ");
// $display("              execution cycles = %7d", total_latency);
// $display("              clock period = %4fns", CYCLE);