NAMESCASESENSITIVE ON ;
MACRO AN2
    CLASS CORE ;
    FOREIGN AN2 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.480 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.000 2.790 2.310 3.190 ;
        RECT  2.030 1.180 2.310 3.300 ;
        RECT  2.000 1.380 2.310 1.780 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.250 1.110 2.650 ;
        RECT  0.790 2.100 1.070 2.740 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 1.650 0.550 2.180 ;
        END
    END I1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.380 2.480 0.380 ;
        RECT  1.340 -0.380 1.740 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.410 4.090 1.810 5.420 ;
        RECT  0.000 4.660 2.480 5.420 ;
        RECT  0.470 4.130 0.870 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.470 3.410 1.760 3.650 ;
        RECT  1.520 1.080 1.760 3.650 ;
        RECT  1.520 2.250 1.790 2.650 ;
        RECT  0.160 1.080 1.760 1.320 ;
    END
END AN2

MACRO AN2B1
    CLASS CORE ;
    FOREIGN AN2B1 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.340 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.340 3.100 2.930 3.340 ;
        RECT  1.600 1.180 3.460 1.420 ;
        RECT  2.650 1.180 2.930 3.340 ;
        END
    END O
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.300 1.070 2.940 ;
        RECT  0.720 2.300 1.070 2.700 ;
        END
    END I1
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.670 2.480 1.950 3.920 ;
        RECT  3.690 2.370 4.170 2.770 ;
        RECT  3.890 2.300 4.170 3.920 ;
        RECT  1.670 3.640 4.170 3.920 ;
        RECT  1.490 2.480 1.950 2.880 ;
        END
    END B1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.330 -0.380 2.730 0.820 ;
        RECT  3.780 -0.380 4.180 1.290 ;
        RECT  0.000 -0.380 4.340 0.380 ;
        RECT  0.880 -0.380 1.280 1.420 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.780 4.160 4.180 5.420 ;
        RECT  0.000 4.660 4.340 5.420 ;
        RECT  0.880 3.910 1.280 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  1.620 4.160 3.460 4.400 ;
        RECT  0.190 3.670 0.480 4.070 ;
        RECT  0.190 1.100 0.430 4.070 ;
        RECT  2.170 1.810 2.410 2.210 ;
        RECT  0.190 1.810 2.410 2.050 ;
        RECT  0.190 1.100 0.480 1.500 ;
    END
END AN2B1

MACRO AN2B1P
    CLASS CORE ;
    FOREIGN AN2B1P 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.960 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.760 2.900 4.170 3.300 ;
        RECT  3.150 1.530 4.800 1.810 ;
        RECT  3.890 1.530 4.170 3.300 ;
        END
    END O
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.100 1.690 2.740 ;
        RECT  1.350 2.100 1.690 2.500 ;
        END
    END I1
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.660 1.070 3.300 ;
        RECT  0.670 2.660 1.070 3.060 ;
        END
    END B1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.780 -0.380 4.180 1.020 ;
        RECT  0.000 -0.380 4.960 0.380 ;
        RECT  1.020 -0.380 1.420 1.130 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.660 4.480 3.060 5.420 ;
        RECT  4.400 4.180 4.800 5.420 ;
        RECT  0.000 4.660 4.960 5.420 ;
        RECT  1.020 3.910 1.420 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  1.850 3.910 2.910 4.150 ;
        RECT  2.670 0.810 2.910 4.150 ;
        RECT  2.670 2.130 3.650 2.530 ;
        RECT  2.510 0.810 2.910 1.210 ;
        RECT  0.190 3.670 0.480 4.070 ;
        RECT  0.190 0.810 0.430 4.070 ;
        RECT  1.930 1.370 2.330 1.690 ;
        RECT  0.190 1.370 2.330 1.610 ;
        RECT  0.190 0.810 0.480 1.610 ;
    END
END AN2B1P

MACRO AN2B1S
    CLASS CORE ;
    FOREIGN AN2B1S 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.100 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 1.070 2.310 2.100 ;
        RECT  2.030 1.820 2.930 2.100 ;
        RECT  2.650 1.820 2.930 3.420 ;
        RECT  2.620 3.020 2.930 3.420 ;
        RECT  1.860 1.070 2.310 1.470 ;
        END
    END O
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 1.610 1.070 2.250 ;
        RECT  0.720 1.610 1.070 2.010 ;
        END
    END I1
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.320 1.700 2.720 ;
        RECT  1.410 2.300 1.690 2.940 ;
        END
    END B1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.550 -0.380 2.940 1.210 ;
        RECT  0.000 -0.380 3.100 0.380 ;
        RECT  1.020 -0.380 1.420 1.230 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 4.660 3.100 5.420 ;
        RECT  1.010 4.480 1.410 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.190 4.000 2.380 4.240 ;
        RECT  2.140 2.480 2.380 4.240 ;
        RECT  0.190 3.830 0.480 4.240 ;
        RECT  0.190 1.070 0.430 4.240 ;
        RECT  2.140 2.480 2.410 2.880 ;
        RECT  0.190 1.070 0.480 1.470 ;
    END
END AN2B1S

MACRO AN2B1T
    CLASS CORE ;
    FOREIGN AN2B1T 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.580 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.750 1.490 5.310 3.280 ;
        RECT  3.610 2.880 5.310 3.280 ;
        RECT  3.610 1.490 5.310 1.890 ;
        END
    END O
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.200 2.630 2.600 ;
        RECT  2.030 2.200 2.310 2.840 ;
        END
    END I1
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.450 1.070 3.400 ;
        RECT  0.740 2.450 1.070 2.850 ;
        END
    END B1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.740 -0.380 3.140 0.560 ;
        RECT  4.260 -0.380 4.660 1.120 ;
        RECT  0.000 -0.380 5.580 0.380 ;
        RECT  0.380 -0.380 0.780 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.910 4.260 3.310 5.420 ;
        RECT  4.260 4.180 4.660 5.420 ;
        RECT  0.000 4.660 5.580 5.420 ;
        RECT  1.400 3.750 1.800 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.120 3.780 3.370 4.020 ;
        RECT  3.130 0.890 3.370 4.020 ;
        RECT  3.130 2.170 3.510 2.570 ;
        RECT  1.400 0.890 3.370 1.130 ;
        RECT  0.240 1.370 0.480 3.390 ;
        RECT  1.430 1.370 1.670 2.310 ;
        RECT  0.240 1.370 1.670 1.610 ;
    END
END AN2B1T

MACRO AN2P
    CLASS CORE ;
    FOREIGN AN2P 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.720 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.520 2.790 2.930 3.190 ;
        RECT  2.650 1.180 2.930 3.300 ;
        RECT  2.520 1.320 2.930 1.720 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.100 1.690 2.740 ;
        RECT  1.360 2.250 1.690 2.650 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 1.540 0.530 1.940 ;
        RECT  0.170 1.540 0.450 2.180 ;
        END
    END I1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.160 -0.380 3.560 0.780 ;
        RECT  0.000 -0.380 3.720 0.380 ;
        RECT  1.670 -0.380 2.070 0.780 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.670 4.260 2.070 5.420 ;
        RECT  3.160 4.260 3.560 5.420 ;
        RECT  0.000 4.660 3.720 5.420 ;
        RECT  0.160 3.780 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.880 3.780 2.280 4.020 ;
        RECT  2.040 1.020 2.280 4.020 ;
        RECT  0.160 1.020 2.280 1.260 ;
    END
END AN2P

MACRO AN2S
    CLASS CORE ;
    FOREIGN AN2S 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.480 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 1.300 2.310 3.400 ;
        RECT  2.000 3.000 2.310 3.400 ;
        RECT  2.000 1.300 2.310 1.700 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.540 1.070 3.300 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 1.840 0.490 2.240 ;
        RECT  0.170 1.740 0.450 2.380 ;
        END
    END I1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.380 2.480 0.380 ;
        RECT  0.900 -0.380 1.300 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.780 4.100 2.180 5.420 ;
        RECT  0.000 4.660 2.480 5.420 ;
        RECT  0.450 4.480 0.850 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.450 3.540 1.760 3.780 ;
        RECT  1.520 0.800 1.760 3.780 ;
        RECT  1.520 2.140 1.770 2.540 ;
        RECT  0.320 0.800 1.760 1.040 ;
        RECT  0.160 0.620 0.560 0.860 ;
    END
END AN2S

MACRO AN2T
    CLASS CORE ;
    FOREIGN AN2T 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.340 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.510 1.490 4.070 3.280 ;
        RECT  2.480 2.880 4.070 3.280 ;
        RECT  2.480 1.490 4.070 1.890 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.530 1.690 3.300 ;
        RECT  1.190 2.530 1.690 2.930 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.100 0.530 2.500 ;
        RECT  0.170 1.740 0.450 2.500 ;
        END
    END I1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.020 -0.380 3.420 1.120 ;
        RECT  0.000 -0.380 4.340 0.380 ;
        RECT  1.540 -0.380 1.940 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.670 4.260 2.070 5.420 ;
        RECT  3.020 4.180 3.420 5.420 ;
        RECT  0.000 4.660 4.340 5.420 ;
        RECT  0.160 3.910 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.880 3.780 2.240 4.020 ;
        RECT  2.000 0.890 2.240 4.020 ;
        RECT  2.000 2.170 2.270 2.570 ;
        RECT  0.160 0.890 2.240 1.130 ;
    END
END AN2T

MACRO AN3
    CLASS CORE ;
    FOREIGN AN3 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.720 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.240 2.790 3.550 3.190 ;
        RECT  3.270 1.180 3.550 3.300 ;
        RECT  3.240 1.490 3.550 1.890 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 1.540 1.690 2.180 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.300 0.530 2.700 ;
        RECT  0.170 2.300 0.450 2.940 ;
        END
    END I1
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.300 2.310 2.940 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.380 3.720 0.380 ;
        RECT  2.370 -0.380 2.770 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.190 4.480 2.590 5.420 ;
        RECT  0.000 4.660 3.720 5.420 ;
        RECT  0.920 4.130 1.320 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.160 3.370 2.910 3.610 ;
        RECT  2.670 0.900 2.910 3.610 ;
        RECT  2.670 2.140 3.030 2.540 ;
        RECT  0.160 0.900 2.910 1.140 ;
        RECT  0.160 0.890 0.560 1.140 ;
    END
END AN3

MACRO AN3B1
    CLASS CORE ;
    FOREIGN AN3B1 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.960 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.480 2.790 4.790 3.190 ;
        RECT  4.510 1.180 4.790 3.300 ;
        RECT  4.480 1.490 4.790 1.890 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 1.640 1.690 2.280 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.840 2.310 3.480 ;
        END
    END I1
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.840 1.070 3.480 ;
        RECT  0.670 2.840 1.070 3.240 ;
        END
    END B1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.610 -0.380 4.010 0.560 ;
        RECT  0.000 -0.380 4.960 0.380 ;
        RECT  0.820 -0.380 1.220 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.130 4.480 2.530 5.420 ;
        RECT  3.680 4.260 4.080 5.420 ;
        RECT  0.000 4.660 4.960 5.420 ;
        RECT  0.950 4.480 1.350 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  1.540 3.720 4.150 3.960 ;
        RECT  3.910 1.020 4.150 3.960 ;
        RECT  3.030 1.020 4.150 1.260 ;
        RECT  3.030 0.860 3.270 1.260 ;
        RECT  0.190 3.570 0.480 3.970 ;
        RECT  0.190 0.940 0.430 3.970 ;
        RECT  2.550 1.500 3.030 1.740 ;
        RECT  2.550 0.940 2.790 1.740 ;
        RECT  0.160 0.940 2.790 1.180 ;
    END
END AN3B1

MACRO AN3B1P
    CLASS CORE ;
    FOREIGN AN3B1P 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.580 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.450 2.790 4.790 3.190 ;
        RECT  4.510 1.180 4.790 3.300 ;
        RECT  4.450 1.320 4.790 1.720 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 1.640 1.690 2.280 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.820 2.310 3.460 ;
        END
    END I1
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.820 1.070 3.460 ;
        RECT  0.670 2.820 1.070 3.220 ;
        END
    END B1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.710 -0.380 4.110 0.860 ;
        RECT  5.020 -0.380 5.420 0.860 ;
        RECT  0.000 -0.380 5.580 0.380 ;
        RECT  0.820 -0.380 1.220 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.200 4.480 2.600 5.420 ;
        RECT  3.710 4.180 4.110 5.420 ;
        RECT  5.020 4.180 5.420 5.420 ;
        RECT  0.000 4.660 5.580 5.420 ;
        RECT  1.020 4.480 1.420 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  1.610 3.700 4.150 3.940 ;
        RECT  3.910 1.100 4.150 3.940 ;
        RECT  3.070 1.100 4.150 1.340 ;
        RECT  3.070 0.940 3.310 1.340 ;
        RECT  0.190 3.580 0.480 3.980 ;
        RECT  0.190 1.020 0.430 3.980 ;
        RECT  2.590 1.580 3.340 1.820 ;
        RECT  2.590 1.020 2.830 1.820 ;
        RECT  0.160 1.020 2.830 1.260 ;
    END
END AN3B1P

MACRO AN3B1S
    CLASS CORE ;
    FOREIGN AN3B1S 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.960 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.510 1.060 4.790 3.710 ;
        RECT  4.480 3.310 4.790 3.710 ;
        RECT  4.480 1.060 4.790 1.460 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 1.540 1.690 2.180 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.300 2.310 2.940 ;
        END
    END I1
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.670 2.540 1.070 2.940 ;
        RECT  0.790 2.300 1.070 2.940 ;
        END
    END B1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.790 -0.380 4.190 0.560 ;
        RECT  0.000 -0.380 4.960 0.380 ;
        RECT  0.820 -0.380 1.220 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.610 4.480 2.010 5.420 ;
        RECT  2.270 4.480 2.670 5.420 ;
        RECT  3.610 4.480 4.010 5.420 ;
        RECT  0.000 4.660 4.960 5.420 ;
        RECT  0.950 4.480 1.350 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  1.540 3.330 4.150 3.570 ;
        RECT  3.910 1.020 4.150 3.570 ;
        RECT  3.150 1.020 4.150 1.260 ;
        RECT  3.150 0.860 3.390 1.260 ;
        RECT  0.190 3.250 0.480 3.650 ;
        RECT  0.190 0.800 0.430 3.650 ;
        RECT  2.670 1.500 3.070 1.740 ;
        RECT  2.670 0.800 2.910 1.740 ;
        RECT  0.160 0.940 0.560 1.180 ;
        RECT  0.190 0.800 2.910 1.040 ;
    END
END AN3B1S

MACRO AN3B1T
    CLASS CORE ;
    FOREIGN AN3B1T 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.200 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.350 2.870 4.590 3.270 ;
        RECT  5.130 1.400 5.410 3.110 ;
        RECT  4.350 1.400 6.040 1.640 ;
        RECT  4.350 2.870 6.040 3.110 ;
        RECT  4.350 1.240 4.590 1.640 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 1.880 1.690 2.750 ;
        RECT  1.350 1.880 1.690 2.280 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.220 2.310 2.860 ;
        END
    END I1
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.220 1.070 2.860 ;
        RECT  0.670 2.220 1.070 2.620 ;
        END
    END B1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.640 -0.380 4.040 0.860 ;
        RECT  5.020 -0.380 5.420 0.860 ;
        RECT  0.000 -0.380 6.200 0.380 ;
        RECT  0.750 -0.380 1.150 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.130 4.480 2.530 5.420 ;
        RECT  3.640 4.180 4.040 5.420 ;
        RECT  5.020 4.180 5.420 5.420 ;
        RECT  0.000 4.660 6.200 5.420 ;
        RECT  0.750 4.480 1.150 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  1.540 3.440 4.080 3.680 ;
        RECT  3.840 1.100 4.080 3.680 ;
        RECT  3.000 1.100 4.080 1.340 ;
        RECT  3.000 0.940 3.240 1.340 ;
        RECT  0.190 3.020 0.480 3.420 ;
        RECT  0.190 1.220 0.430 3.420 ;
        RECT  2.500 1.820 3.090 2.060 ;
        RECT  2.500 1.220 2.740 2.060 ;
        RECT  0.160 1.280 0.560 1.520 ;
        RECT  0.190 1.220 2.740 1.460 ;
    END
END AN3B1T

MACRO AN3B2
    CLASS CORE ;
    FOREIGN AN3B2 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.580 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.100 2.790 5.410 3.190 ;
        RECT  5.130 1.180 5.410 3.300 ;
        RECT  5.100 1.490 5.410 1.890 ;
        END
    END O
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.220 1.540 1.690 1.940 ;
        RECT  1.410 0.960 1.690 1.940 ;
        END
    END I1
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.760 1.070 3.400 ;
        RECT  0.710 2.760 1.070 3.160 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.890 2.100 4.170 2.740 ;
        END
    END B1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.130 -0.380 4.530 0.560 ;
        RECT  0.000 -0.380 5.580 0.380 ;
        RECT  0.820 -0.380 1.220 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.230 4.480 2.630 5.420 ;
        RECT  4.250 4.480 4.650 5.420 ;
        RECT  0.000 4.660 5.580 5.420 ;
        RECT  0.750 4.480 1.150 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  1.620 4.000 4.770 4.240 ;
        RECT  4.530 0.800 4.770 4.240 ;
        RECT  3.000 3.640 3.240 4.240 ;
        RECT  1.620 3.640 1.860 4.240 ;
        RECT  4.530 2.140 4.870 2.540 ;
        RECT  2.650 0.800 4.770 1.040 ;
        RECT  3.050 1.490 3.290 3.190 ;
        RECT  2.950 2.030 3.290 2.430 ;
        RECT  3.050 1.490 3.340 1.890 ;
        RECT  0.190 3.580 0.480 3.980 ;
        RECT  0.190 0.860 0.430 3.980 ;
        RECT  0.190 2.280 2.130 2.520 ;
        RECT  0.190 0.860 0.480 1.260 ;
    END
END AN3B2

MACRO AN3B2P
    CLASS CORE ;
    FOREIGN AN3B2P 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.200 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.100 2.790 5.410 3.190 ;
        RECT  5.130 1.180 5.410 3.300 ;
        RECT  5.100 1.490 5.410 1.890 ;
        END
    END O
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.310 1.540 1.690 1.940 ;
        RECT  1.410 1.180 1.690 1.940 ;
        END
    END I1
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.760 1.070 3.400 ;
        RECT  0.710 2.760 1.070 3.160 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.890 2.100 4.170 2.740 ;
        END
    END B1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.130 -0.380 4.530 0.560 ;
        RECT  5.640 -0.380 6.040 1.070 ;
        RECT  0.000 -0.380 6.200 0.380 ;
        RECT  0.820 -0.380 1.220 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.330 4.480 2.730 5.420 ;
        RECT  4.400 4.220 4.800 5.420 ;
        RECT  5.640 4.220 6.040 5.420 ;
        RECT  0.000 4.660 6.200 5.420 ;
        RECT  0.750 4.480 1.150 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  1.540 3.660 4.770 3.900 ;
        RECT  4.530 0.800 4.770 3.900 ;
        RECT  4.530 2.140 4.870 2.540 ;
        RECT  2.670 0.800 4.770 1.040 ;
        RECT  3.290 1.490 3.530 3.190 ;
        RECT  3.050 2.100 3.530 2.500 ;
        RECT  0.190 3.580 0.480 3.980 ;
        RECT  0.190 0.930 0.430 3.980 ;
        RECT  0.190 2.280 2.310 2.520 ;
        RECT  0.190 0.930 0.480 1.330 ;
    END
END AN3B2P

MACRO AN3B2S
    CLASS CORE ;
    FOREIGN AN3B2S 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.720 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.270 1.120 3.550 3.300 ;
        RECT  3.240 2.900 3.550 3.300 ;
        RECT  1.600 1.140 3.560 1.380 ;
        RECT  1.600 1.120 3.550 1.400 ;
        END
    END O
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 1.690 1.070 2.330 ;
        RECT  0.720 1.690 1.070 2.090 ;
        END
    END I1
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.100 1.690 2.740 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 1.690 2.350 2.090 ;
        RECT  2.030 1.690 2.310 2.330 ;
        END
    END B1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.370 -0.380 2.770 0.560 ;
        RECT  0.000 -0.380 3.720 0.380 ;
        RECT  0.880 -0.380 1.280 1.380 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 4.660 3.720 5.420 ;
        RECT  1.040 4.260 1.440 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.190 3.780 3.000 4.020 ;
        RECT  2.760 2.250 3.000 4.020 ;
        RECT  0.190 3.620 0.480 4.020 ;
        RECT  0.190 1.060 0.430 4.020 ;
        RECT  2.760 2.250 3.030 2.650 ;
        RECT  0.190 1.060 0.480 1.460 ;
    END
END AN3B2S

MACRO AN3B2T
    CLASS CORE ;
    FOREIGN AN3B2T 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.820 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.100 2.870 5.340 3.270 ;
        RECT  5.750 1.570 6.030 3.110 ;
        RECT  5.100 1.570 6.660 1.810 ;
        RECT  5.100 2.870 6.660 3.110 ;
        RECT  5.100 1.410 5.340 1.810 ;
        END
    END O
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.310 1.540 1.690 1.940 ;
        RECT  1.410 1.180 1.690 1.940 ;
        END
    END I1
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.660 1.070 3.400 ;
        RECT  0.710 2.660 1.070 3.060 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.890 1.880 4.170 2.520 ;
        END
    END B1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.130 -0.380 4.530 0.560 ;
        RECT  5.640 -0.380 6.040 1.070 ;
        RECT  0.000 -0.380 6.820 0.380 ;
        RECT  0.820 -0.380 1.220 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.330 4.480 2.730 5.420 ;
        RECT  4.400 4.220 4.800 5.420 ;
        RECT  5.640 4.220 6.040 5.420 ;
        RECT  0.000 4.660 6.820 5.420 ;
        RECT  0.750 4.480 1.150 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  1.540 3.660 4.770 3.900 ;
        RECT  4.530 0.820 4.770 3.900 ;
        RECT  4.530 2.140 4.870 2.540 ;
        RECT  2.670 0.820 4.770 1.060 ;
        RECT  3.290 2.870 4.010 3.110 ;
        RECT  3.290 1.490 3.530 3.110 ;
        RECT  3.050 2.100 3.530 2.500 ;
        RECT  0.190 3.580 0.480 3.980 ;
        RECT  0.190 0.930 0.430 3.980 ;
        RECT  0.190 2.180 2.310 2.420 ;
        RECT  0.190 0.930 0.480 1.330 ;
    END
END AN3B2T

MACRO AN3P
    CLASS CORE ;
    FOREIGN AN3P 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.340 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.140 2.790 3.550 3.190 ;
        RECT  3.270 1.180 3.550 3.300 ;
        RECT  3.140 1.490 3.550 1.890 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.300 1.690 2.940 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 1.540 0.530 1.940 ;
        RECT  0.170 1.540 0.450 2.180 ;
        END
    END I1
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 1.540 2.310 2.180 ;
        RECT  1.980 1.540 2.310 1.940 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.780 -0.380 4.180 0.950 ;
        RECT  0.000 -0.380 4.340 0.380 ;
        RECT  2.150 -0.380 2.550 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.330 4.260 2.730 5.420 ;
        RECT  3.780 4.260 4.180 5.420 ;
        RECT  0.000 4.660 4.340 5.420 ;
        RECT  0.850 4.130 1.250 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.160 3.360 2.900 3.600 ;
        RECT  2.660 0.890 2.900 3.600 ;
        RECT  0.160 0.890 2.900 1.130 ;
    END
END AN3P

MACRO AN3S
    CLASS CORE ;
    FOREIGN AN3S 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.720 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.270 0.620 3.550 3.850 ;
        RECT  3.240 3.450 3.550 3.850 ;
        RECT  3.240 0.670 3.550 1.070 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 1.540 1.690 2.180 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.100 0.550 2.500 ;
        RECT  0.170 2.100 0.450 2.740 ;
        END
    END I1
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.100 2.310 2.740 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.380 3.720 0.380 ;
        RECT  2.370 -0.380 2.770 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.370 4.130 2.770 5.420 ;
        RECT  0.000 4.660 3.720 5.420 ;
        RECT  0.920 4.130 1.320 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.160 3.370 2.910 3.610 ;
        RECT  2.670 0.800 2.910 3.610 ;
        RECT  2.670 2.140 3.030 2.540 ;
        RECT  0.160 0.800 0.560 1.130 ;
        RECT  0.160 0.800 2.910 1.040 ;
    END
END AN3S

MACRO AN3T
    CLASS CORE ;
    FOREIGN AN3T 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.960 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.040 2.870 3.280 3.270 ;
        RECT  3.890 1.570 4.170 3.110 ;
        RECT  3.040 1.570 4.800 1.810 ;
        RECT  3.040 2.870 4.800 3.110 ;
        RECT  3.040 1.410 3.280 1.810 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.090 1.690 2.790 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 1.620 0.530 2.020 ;
        RECT  0.170 1.620 0.450 2.260 ;
        END
    END I1
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 1.620 2.310 2.260 ;
        RECT  1.930 1.620 2.310 2.020 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.680 -0.380 4.080 0.950 ;
        RECT  0.000 -0.380 4.960 0.380 ;
        RECT  2.150 -0.380 2.550 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.240 4.260 2.640 5.420 ;
        RECT  3.680 4.260 4.080 5.420 ;
        RECT  0.000 4.660 4.960 5.420 ;
        RECT  0.850 4.130 1.250 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.160 3.360 2.790 3.600 ;
        RECT  2.550 0.890 2.790 3.600 ;
        RECT  2.550 2.140 3.400 2.540 ;
        RECT  0.160 0.890 2.790 1.130 ;
    END
END AN3T

MACRO AN4
    CLASS CORE ;
    FOREIGN AN4 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.200 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.130 1.420 5.410 3.260 ;
        RECT  4.500 2.860 5.410 3.260 ;
        RECT  4.800 1.420 5.410 1.660 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.400 1.260 2.800 ;
        RECT  0.790 2.160 1.070 2.800 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 1.910 0.500 2.310 ;
        RECT  0.170 1.540 0.450 2.310 ;
        END
    END I1
    PIN I4
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.930 1.910 2.310 2.310 ;
        RECT  2.030 1.540 2.310 2.310 ;
        END
    END I4
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 2.160 2.930 2.800 ;
        RECT  2.610 2.260 2.930 2.660 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.910 -0.380 4.310 0.560 ;
        RECT  5.640 -0.380 6.040 0.810 ;
        RECT  0.000 -0.380 6.200 0.380 ;
        RECT  1.450 -0.380 1.850 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.920 4.480 3.320 5.420 ;
        RECT  5.640 4.260 6.040 5.420 ;
        RECT  0.000 4.660 6.200 5.420 ;
        RECT  0.160 4.480 1.740 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.830 4.000 4.770 4.240 ;
        RECT  5.710 2.300 5.950 4.020 ;
        RECT  4.530 3.780 5.950 4.020 ;
        RECT  0.830 3.040 1.070 4.240 ;
        RECT  0.830 3.040 3.410 3.280 ;
        RECT  3.170 0.800 3.410 3.280 ;
        RECT  3.170 2.060 3.530 2.460 ;
        RECT  0.160 0.800 0.560 1.130 ;
        RECT  0.160 0.800 3.410 1.040 ;
        RECT  2.130 3.520 4.260 3.760 ;
        RECT  4.020 1.470 4.260 3.760 ;
        RECT  4.020 2.380 4.590 2.620 ;
        RECT  3.650 1.470 4.260 1.710 ;
        RECT  3.650 1.310 3.890 1.710 ;
    END
END AN4

MACRO AN4B1
    CLASS CORE ;
    FOREIGN AN4B1 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.580 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.830 2.930 4.170 3.330 ;
        RECT  3.890 1.280 4.650 1.560 ;
        RECT  3.890 1.280 4.170 3.330 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.350 1.760 1.690 2.160 ;
        RECT  1.410 1.180 1.690 2.160 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.300 2.310 2.940 ;
        END
    END I1
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.100 1.590 3.550 1.990 ;
        RECT  3.270 0.800 5.410 1.040 ;
        RECT  4.870 2.300 5.410 2.700 ;
        RECT  5.130 0.800 5.410 2.740 ;
        RECT  3.270 0.800 3.550 1.990 ;
        END
    END B1
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.300 0.490 2.700 ;
        RECT  0.170 2.300 0.450 2.940 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.440 -0.380 3.840 0.560 ;
        RECT  5.020 -0.380 5.420 0.560 ;
        RECT  0.000 -0.380 5.580 0.380 ;
        RECT  0.160 -0.380 0.560 0.780 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.190 4.480 2.590 5.420 ;
        RECT  5.020 4.260 5.420 5.420 ;
        RECT  0.000 4.660 5.580 5.420 ;
        RECT  0.830 4.480 1.230 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.160 3.690 2.800 3.930 ;
        RECT  2.560 1.220 2.800 3.930 ;
        RECT  3.410 2.290 3.650 2.690 ;
        RECT  2.560 2.350 3.650 2.590 ;
    END
END AN4B1

MACRO AN4B1P
    CLASS CORE ;
    FOREIGN AN4B1P 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.060 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.840 2.940 6.680 3.220 ;
        RECT  3.320 1.260 7.900 1.540 ;
        RECT  4.510 1.260 4.790 3.220 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 1.540 1.690 2.430 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.300 2.400 2.700 ;
        RECT  2.030 2.300 2.310 2.940 ;
        END
    END I1
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.170 2.380 5.570 2.620 ;
        RECT  5.330 1.790 7.890 2.030 ;
        RECT  7.410 1.790 7.890 2.700 ;
        RECT  7.610 1.790 7.890 2.740 ;
        RECT  5.330 1.790 5.570 2.620 ;
        END
    END B1
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.300 0.490 2.700 ;
        RECT  0.170 2.300 0.450 2.940 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.830 -0.380 4.230 0.560 ;
        RECT  5.410 -0.380 5.810 0.560 ;
        RECT  6.710 -0.380 7.110 0.560 ;
        RECT  0.000 -0.380 8.060 0.380 ;
        RECT  0.160 -0.380 0.560 0.780 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.640 4.260 3.040 5.420 ;
        RECT  5.060 4.260 5.460 5.420 ;
        RECT  7.500 4.260 7.900 5.420 ;
        RECT  0.000 4.660 8.060 5.420 ;
        RECT  0.950 4.480 1.350 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.160 3.780 3.080 4.020 ;
        RECT  2.840 0.620 3.080 4.020 ;
        RECT  6.920 2.380 7.160 3.780 ;
        RECT  2.840 3.540 7.160 3.780 ;
        RECT  6.330 2.380 7.160 2.620 ;
        RECT  2.840 2.370 4.010 2.610 ;
        RECT  2.390 0.620 3.080 1.020 ;
    END
END AN4B1P

MACRO AN4B1S
    CLASS CORE ;
    FOREIGN AN4B1S 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.340 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.860 0.640 4.170 1.040 ;
        RECT  2.130 0.800 4.170 1.040 ;
        RECT  3.860 3.220 4.170 3.620 ;
        RECT  3.890 0.640 4.170 3.860 ;
        RECT  2.130 0.720 2.530 1.040 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 0.920 1.690 1.620 ;
        RECT  1.330 0.920 1.690 1.320 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.100 2.310 2.740 ;
        RECT  2.010 2.100 2.310 2.500 ;
        END
    END I1
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 2.680 3.050 3.080 ;
        RECT  2.650 2.680 2.930 3.300 ;
        END
    END B1
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 2.100 0.550 2.500 ;
        RECT  0.170 2.100 0.450 2.740 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.990 -0.380 3.390 0.560 ;
        RECT  0.000 -0.380 4.340 0.380 ;
        RECT  0.240 -0.380 0.480 1.190 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.370 4.480 2.770 5.420 ;
        RECT  0.000 4.660 4.340 5.420 ;
        RECT  0.720 4.480 1.120 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.160 3.650 3.530 3.890 ;
        RECT  3.290 1.280 3.530 3.890 ;
        RECT  2.450 1.280 2.690 1.860 ;
        RECT  3.290 1.280 3.650 1.680 ;
        RECT  2.450 1.280 3.650 1.520 ;
    END
END AN4B1S

MACRO AN4B1T
    CLASS CORE ;
    FOREIGN AN4B1T 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.540 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.860 2.960 4.140 3.340 ;
        RECT  8.870 1.350 9.110 3.200 ;
        RECT  3.860 2.960 9.110 3.200 ;
        RECT  3.850 1.350 10.380 1.590 ;
        RECT  3.860 2.940 4.100 3.340 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.370 2.250 1.690 2.650 ;
        RECT  1.410 1.910 1.690 2.650 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 2.250 2.330 2.650 ;
        RECT  2.030 2.160 2.310 2.800 ;
        END
    END I1
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 2.250 3.080 2.650 ;
        RECT  2.650 3.580 4.720 3.820 ;
        RECT  4.480 3.540 9.730 3.780 ;
        RECT  9.490 2.250 9.730 3.780 ;
        RECT  9.490 2.250 9.970 2.650 ;
        RECT  2.650 2.160 2.930 3.820 ;
        END
    END B1
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.790 2.100 1.070 2.740 ;
        RECT  0.690 2.250 1.070 2.650 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.570 -0.380 4.970 1.030 ;
        RECT  6.010 -0.380 6.410 1.030 ;
        RECT  7.820 -0.380 8.220 1.030 ;
        RECT  9.260 -0.380 9.660 1.030 ;
        RECT  0.000 -0.380 10.540 0.380 ;
        RECT  0.160 -0.380 0.560 0.800 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.400 4.260 2.800 5.420 ;
        RECT  4.960 4.260 5.360 5.420 ;
        RECT  7.400 4.260 7.800 5.420 ;
        RECT  9.890 4.260 10.290 5.420 ;
        RECT  0.000 4.660 10.540 5.420 ;
        RECT  0.880 3.910 1.280 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.160 3.430 2.010 3.670 ;
        RECT  0.160 1.150 0.400 3.670 ;
        RECT  8.390 2.280 8.630 2.680 ;
        RECT  3.320 2.330 8.630 2.570 ;
        RECT  3.320 1.150 3.560 2.570 ;
        RECT  3.210 1.150 3.560 1.670 ;
        RECT  0.160 1.150 3.560 1.390 ;
    END
END AN4B1T

MACRO AN4P
    CLASS CORE ;
    FOREIGN AN4P 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.680 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.490 2.940 4.790 3.340 ;
        RECT  4.110 0.800 4.770 1.040 ;
        RECT  4.530 0.800 4.770 1.540 ;
        RECT  4.510 2.940 4.790 3.860 ;
        RECT  7.610 1.260 7.890 3.220 ;
        RECT  4.490 2.940 7.890 3.220 ;
        RECT  4.530 1.260 8.520 1.540 ;
        RECT  3.800 0.620 4.350 0.860 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.100 1.690 2.740 ;
        RECT  1.310 2.250 1.690 2.650 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 1.880 0.500 2.280 ;
        RECT  0.170 1.540 0.450 2.280 ;
        END
    END I1
    PIN I4
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.990 1.880 2.310 2.280 ;
        RECT  2.030 1.540 2.310 2.280 ;
        END
    END I4
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 2.250 2.950 2.650 ;
        RECT  2.650 2.160 2.930 2.800 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  4.590 -0.380 4.990 0.560 ;
        RECT  6.030 -0.380 6.430 0.560 ;
        RECT  7.330 -0.380 7.730 0.560 ;
        RECT  0.000 -0.380 8.680 0.380 ;
        RECT  1.550 -0.380 1.950 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.930 4.480 3.330 5.420 ;
        RECT  5.590 4.260 5.990 5.420 ;
        RECT  8.030 4.260 8.430 5.420 ;
        RECT  0.000 4.660 8.680 5.420 ;
        RECT  0.160 4.480 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.910 4.160 5.350 4.400 ;
        RECT  5.110 3.540 5.350 4.400 ;
        RECT  1.590 4.000 4.150 4.240 ;
        RECT  1.590 3.040 1.830 4.240 ;
        RECT  5.110 3.540 8.370 3.780 ;
        RECT  8.130 2.300 8.370 3.780 ;
        RECT  0.750 3.040 3.530 3.280 ;
        RECT  3.290 0.800 3.530 3.280 ;
        RECT  3.290 2.030 3.670 2.430 ;
        RECT  0.160 0.800 3.530 1.040 ;
        RECT  2.140 3.520 4.150 3.760 ;
        RECT  3.910 1.340 4.150 3.760 ;
        RECT  3.910 2.380 7.260 2.620 ;
        RECT  3.830 1.340 4.150 1.740 ;
    END
END AN4P

MACRO AN4S
    CLASS CORE ;
    FOREIGN AN4S 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.960 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.350 3.350 4.790 3.750 ;
        RECT  4.510 0.850 4.790 3.860 ;
        RECT  3.810 0.850 4.790 1.130 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.970 2.360 1.210 2.760 ;
        RECT  0.790 2.100 1.070 2.740 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 1.540 0.500 1.940 ;
        RECT  0.170 1.540 0.450 2.180 ;
        END
    END I1
    PIN I4
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.930 2.860 2.390 3.300 ;
        END
    END I4
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.630 2.860 3.050 3.300 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.020 -0.380 3.420 0.560 ;
        RECT  0.000 -0.380 4.960 0.380 ;
        RECT  1.410 -0.380 1.810 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.950 4.480 3.350 5.420 ;
        RECT  0.000 4.660 4.960 5.420 ;
        RECT  0.160 4.480 1.740 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  2.130 3.940 4.110 4.180 ;
        RECT  3.870 1.370 4.110 4.180 ;
        RECT  3.870 2.300 4.270 2.700 ;
        RECT  2.500 1.370 4.110 1.610 ;
        RECT  0.750 3.650 1.690 3.890 ;
        RECT  1.450 0.890 1.690 3.890 ;
        RECT  1.450 1.850 3.630 2.090 ;
        RECT  0.160 0.890 1.690 1.130 ;
    END
END AN4S

MACRO AN4T
    CLASS CORE ;
    FOREIGN AN4T 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.160 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.520 2.960 4.760 3.860 ;
        RECT  9.490 1.350 9.730 3.200 ;
        RECT  4.480 2.960 9.730 3.200 ;
        RECT  4.470 1.350 11.000 1.590 ;
        RECT  4.480 2.940 4.720 3.340 ;
        END
    END O
    PIN I2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.100 1.690 2.740 ;
        RECT  1.310 2.250 1.690 2.650 ;
        END
    END I2
    PIN I1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 1.880 0.500 2.280 ;
        RECT  0.170 1.540 0.450 2.280 ;
        END
    END I1
    PIN I4
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.990 1.880 2.310 2.280 ;
        RECT  2.030 1.540 2.310 2.280 ;
        END
    END I4
    PIN I3
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 2.250 2.950 2.650 ;
        RECT  2.650 2.160 2.930 2.800 ;
        END
    END I3
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  5.190 -0.380 5.590 1.030 ;
        RECT  6.630 -0.380 7.030 1.030 ;
        RECT  8.440 -0.380 8.840 1.030 ;
        RECT  9.880 -0.380 10.280 1.030 ;
        RECT  0.000 -0.380 11.160 0.380 ;
        RECT  1.550 -0.380 1.950 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.930 4.480 3.330 5.420 ;
        RECT  5.580 4.260 5.980 5.420 ;
        RECT  8.020 4.260 8.420 5.420 ;
        RECT  10.510 4.260 10.910 5.420 ;
        RECT  0.000 4.660 11.160 5.420 ;
        RECT  0.160 4.480 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.900 4.160 5.340 4.400 ;
        RECT  5.100 3.540 5.340 4.400 ;
        RECT  1.590 4.000 4.140 4.240 ;
        RECT  1.590 3.040 1.830 4.240 ;
        RECT  5.100 3.540 10.660 3.780 ;
        RECT  10.420 2.250 10.660 3.780 ;
        RECT  0.750 3.040 3.530 3.280 ;
        RECT  3.290 0.800 3.530 3.280 ;
        RECT  10.360 2.250 10.660 2.650 ;
        RECT  3.290 2.030 3.670 2.430 ;
        RECT  0.160 0.800 3.530 1.040 ;
        RECT  2.130 3.520 4.180 3.760 ;
        RECT  3.940 1.270 4.180 3.760 ;
        RECT  9.010 2.280 9.250 2.680 ;
        RECT  3.940 2.330 9.250 2.570 ;
        RECT  3.830 1.270 4.180 1.670 ;
    END
END AN4T

MACRO ANTENNA
    CLASS CORE ANTENNACELL ;
    FOREIGN ANTENNA 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.240 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 1.180 1.070 1.620 ;
        END
    END A
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 -0.380 1.240 0.380 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 4.660 1.240 5.420 ;
        END
    END VCC
END ANTENNA

MACRO AO112
    CLASS CORE ;
    FOREIGN AO112 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.960 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 1.300 0.480 1.700 ;
        RECT  0.170 2.790 0.480 3.190 ;
        RECT  0.170 1.300 0.450 3.190 ;
        END
    END O
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.270 2.240 3.650 2.640 ;
        RECT  3.270 2.160 3.550 2.740 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.510 1.530 4.790 2.180 ;
        RECT  4.470 1.530 4.790 1.930 ;
        END
    END A1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.160 1.690 2.810 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 1.570 2.360 1.970 ;
        RECT  2.030 1.530 2.310 2.180 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.460 -0.380 3.860 0.560 ;
        RECT  0.000 -0.380 4.960 0.380 ;
        RECT  1.050 -0.380 1.450 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.450 4.480 2.850 5.420 ;
        RECT  0.000 4.660 4.960 5.420 ;
        RECT  0.740 4.480 1.140 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.910 3.910 4.800 4.150 ;
        RECT  3.910 0.890 4.150 4.150 ;
        RECT  0.700 2.150 1.050 2.550 ;
        RECT  0.810 0.890 1.050 2.550 ;
        RECT  0.810 0.890 4.790 1.130 ;
        RECT  1.530 3.910 3.590 4.150 ;
    END
END AO112

MACRO AO112P
    CLASS CORE ;
    FOREIGN AO112P 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.580 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.960 1.220 1.200 1.620 ;
        RECT  0.170 1.380 1.200 1.620 ;
        RECT  0.170 2.870 1.280 3.110 ;
        RECT  0.170 1.380 0.450 3.110 ;
        END
    END O
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.890 2.240 4.280 2.640 ;
        RECT  3.890 1.950 4.170 2.880 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.130 1.950 5.410 2.880 ;
        RECT  5.090 2.250 5.410 2.650 ;
        END
    END A1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 1.950 2.310 2.890 ;
        RECT  1.950 2.250 2.310 2.650 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 1.950 2.930 2.890 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 -0.380 2.000 0.950 ;
        RECT  4.230 -0.380 4.630 1.230 ;
        RECT  0.000 -0.380 5.580 0.380 ;
        RECT  0.160 -0.380 0.560 0.950 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  1.600 4.170 2.000 5.420 ;
        RECT  3.050 3.930 3.450 5.420 ;
        RECT  0.000 4.660 5.580 5.420 ;
        RECT  0.160 4.170 0.560 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  4.530 3.910 5.420 4.150 ;
        RECT  4.530 1.470 4.770 4.150 ;
        RECT  1.190 2.150 1.680 2.550 ;
        RECT  1.440 1.470 1.680 2.550 ;
        RECT  1.440 1.470 5.420 1.710 ;
        RECT  2.330 3.450 4.030 3.690 ;
        RECT  3.640 3.210 4.040 3.450 ;
    END
END AO112P

MACRO AO112S
    CLASS CORE ;
    FOREIGN AO112S 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.960 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 0.810 0.480 1.210 ;
        RECT  0.170 3.330 0.510 3.730 ;
        RECT  0.170 0.810 0.450 3.730 ;
        END
    END O
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.270 2.790 3.560 3.190 ;
        RECT  3.270 2.720 3.550 3.370 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.510 2.090 4.790 2.740 ;
        RECT  4.410 2.180 4.790 2.580 ;
        END
    END A1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.720 1.690 3.370 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.030 1.640 2.310 2.290 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.460 -0.380 3.860 0.570 ;
        RECT  0.000 -0.380 4.960 0.380 ;
        RECT  1.040 -0.380 1.440 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.470 4.480 2.870 5.420 ;
        RECT  0.000 4.660 4.960 5.420 ;
        RECT  0.890 4.480 1.290 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  3.910 3.870 4.800 4.110 ;
        RECT  3.910 0.890 4.150 4.110 ;
        RECT  0.720 1.350 1.050 1.750 ;
        RECT  0.810 0.890 1.050 1.750 ;
        RECT  0.810 0.890 4.800 1.130 ;
        RECT  1.680 3.870 3.590 4.110 ;
    END
END AO112S

MACRO AO112T
    CLASS CORE ;
    FOREIGN AO112T 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.200 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.680 1.220 1.920 1.620 ;
        RECT  0.160 1.380 1.920 1.620 ;
        RECT  0.160 2.870 2.000 3.110 ;
        RECT  0.790 1.380 1.070 3.110 ;
        END
    END O
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  4.510 2.240 4.900 2.640 ;
        RECT  4.510 1.940 4.790 2.880 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  5.750 1.950 6.030 2.880 ;
        RECT  5.710 2.250 6.030 2.650 ;
        END
    END A1
    PIN C2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.650 1.950 2.930 2.890 ;
        RECT  2.640 2.250 2.930 2.650 ;
        END
    END C2
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.270 2.250 3.620 2.650 ;
        RECT  3.270 1.950 3.550 2.890 ;
        END
    END C1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.320 -0.380 2.720 0.950 ;
        RECT  4.850 -0.380 5.250 1.170 ;
        RECT  0.000 -0.380 6.200 0.380 ;
        RECT  0.880 -0.380 1.280 0.950 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.320 4.170 2.720 5.420 ;
        RECT  3.770 3.930 4.170 5.420 ;
        RECT  0.000 4.660 6.200 5.420 ;
        RECT  0.880 4.170 1.280 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  5.150 3.910 6.040 4.150 ;
        RECT  5.150 1.410 5.390 4.150 ;
        RECT  1.910 2.150 2.400 2.550 ;
        RECT  2.160 1.410 2.400 2.550 ;
        RECT  2.160 1.410 6.040 1.650 ;
        RECT  3.050 3.450 4.750 3.690 ;
        RECT  4.340 3.210 4.740 3.690 ;
    END
END AO112T

MACRO AO12
    CLASS CORE ;
    FOREIGN AO12 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.720 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.270 0.620 3.550 3.290 ;
        RECT  3.170 2.890 3.550 3.290 ;
        RECT  3.240 1.260 3.550 1.660 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 1.510 0.490 1.910 ;
        RECT  0.170 1.090 0.450 1.910 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.100 1.690 2.890 ;
        RECT  1.310 2.100 1.690 2.500 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.020 2.120 2.310 2.520 ;
        RECT  2.030 1.730 2.310 2.520 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.240 -0.380 2.640 0.560 ;
        RECT  0.000 -0.380 3.720 0.380 ;
        RECT  0.160 -0.380 0.560 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  0.000 4.660 3.720 5.420 ;
        RECT  2.430 4.250 2.830 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.880 3.420 1.280 3.760 ;
        RECT  0.880 3.420 2.910 3.660 ;
        RECT  2.670 0.890 2.910 3.660 ;
        RECT  2.670 2.150 3.030 2.550 ;
        RECT  1.440 0.890 2.910 1.130 ;
        RECT  0.160 4.000 2.000 4.240 ;
        RECT  1.600 3.900 2.000 4.240 ;
        RECT  0.160 3.770 0.560 4.240 ;
    END
END AO12

MACRO AO12P
    CLASS CORE ;
    FOREIGN AO12P 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.340 BY 5.040 ;
    SYMMETRY x y   ;
    SITE core_5040 ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT  3.270 1.150 3.550 3.260 ;
        RECT  3.170 2.860 3.550 3.260 ;
        RECT  3.140 1.260 3.550 1.660 ;
        END
    END O
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  0.170 1.710 0.490 2.110 ;
        RECT  0.170 1.540 0.450 2.180 ;
        END
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  1.410 2.100 1.690 2.890 ;
        RECT  1.310 2.100 1.690 2.500 ;
        END
    END B1
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT  2.020 2.120 2.310 2.520 ;
        RECT  2.030 1.730 2.310 2.520 ;
        END
    END A1
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  2.240 -0.380 2.640 0.560 ;
        RECT  3.780 -0.380 4.180 0.930 ;
        RECT  0.000 -0.380 4.340 0.380 ;
        RECT  0.160 -0.380 0.560 0.560 ;
        END
    END GND
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        CLASS CORE ;
        LAYER metal1 ;
        RECT  3.780 4.180 4.180 5.420 ;
        RECT  0.000 4.660 4.340 5.420 ;
        RECT  2.430 4.180 2.830 5.420 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        RECT  0.880 3.400 2.800 3.640 ;
        RECT  2.560 0.890 2.800 3.640 ;
        RECT  2.560 2.150 3.030 2.550 ;
        RECT  1.440 0.890 2.800 1.130 ;
        RECT  0.160 3.880 2.000 4.120 ;
    END
END AO12P

MACRO AO12S
    CLASS CORE ;
    FOREIGN AO12S 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.720 BY 5.040 ;
    SYMMETRY