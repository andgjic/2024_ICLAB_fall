/**************************************************************************/
// Copyright (c) 2024, OASIS Lab
// MODULE: PATTERN
// FILE NAME: PATTERN.v
// VERSRION: 1.0
// DATE: August 15, 2024
// AUTHOR: Yu-Hsuan Hsu, NYCU IEE
// DESCRIPTION: ICLAB2024FALL / LAB3 / PATTERN
// MODIFICATION HISTORY:
// Date                 Description
// 
/**************************************************************************/

`ifdef RTL
    `define CYCLE_TIME 40.0
`endif
`ifdef GATE
    `define CYCLE_TIME 40.0
`endif

module PATTERN(
	//OUTPUT
	rst_n,
	clk,
	in_valid,
	tetrominoes,
	position,
	//INPUT
	tetris_valid,
	score_valid,
	fail,
	score,
	tetris
);


`protected
6N[?]YL,]=2T\O.\Q:-Z<TDE4UUK5A:0Q<F5=H]cJC/Lf-=f/cZ-7)N\-Q#b-CL=
Dd,>c@0P>&@824P8#L+;G?96:O)4?<EJ1eUA<WINV(AK=OKFR.R_a+ANHRO95?^0
fTO#<S@,XSfcY(UEM\dKTZdW.>#NC2Y-@.#B0Z\Ube[UX[R^@FcAZ>DM#g4)=#f,
X#H^7IPRQJ_DaI:2CUO@aKa/EU2aW<9VC/-e/(8STR),(:P+@/AJ5]-KY036Kd0P
,X+NY\8;gcS&+[F8AS0X:]ae^?&P6,A]b-]TYCeIF)]]LFB(8.#<U;-KK$
`endprotected
output reg			rst_n, clk, in_valid;
output reg	[2:0]	tetrominoes;
output reg  [2:0]	position;
input 				tetris_valid, score_valid, fail;
input 		[3:0]	score;
input		[71:0]	tetris;


`protected
bX5Z<eKV^CKZbUEOCP_&8:b:Lf,99Ua^GJIVeCd:JXS)d8gXJD\-+)CL:H+C7K<<
8J80P,>ZVaKT=GUO0JJ\6cF]?)EP=VAbIBKLG8UMZ2ECVVTWb/e:&<^@RB\0Kg/@
7RK2AK:?WgGVU&8,,DM>)[BYe][S<[?YOJ0,Ta)4fN6OV4WZD5EF\L@65)&AM1(d
<22=&5,6IdU>#3,QKEeD?N5@0J2b,SPSb5WH3cQRTO9G]_<R-@A<8)bO5:d0Y0&&
CTUL?fT):\SBNIGgE4@-;\#[R99_=Z@@._WdR)44HLH=a8,Y>H@DB:,T)ggV/T.0
VD26-8?/I.P84LeKX0#61L@c,(W/U=FJ9Y\d)e\F?P(5^G5Q?3H)eM7HaeDP8(YK
R71,,;dYP4Ead:?eNIaD:87:N?3+<=?J[.EPG14J3gE#YfT5LZMA,;(5VbBB\\-<
@&RASeQY4FU?TW0[MAATHaVc=gQ;@SZbPHafEZ4HNS#XI>gUWEBL4<#0YJF;MJJ<
?8R.5cCbd32&#)V8S75fV_7B.0;0f:N1_+XXHJ3(?MX6f5TXBRge(9S8H[^:a7=(
G+_&NE3O;R>ZL2?gf#8Y/0/+T/AD_/cUVF@b>+SfHM:_H8Q^#V^Wc[-F:WJWA+fQ
R]Z;,gJCPRSW927#?2b[@NaKW#8M[Sc;G9+>FP.LV^7ad+RNKM/gG?G,=fYOR>IQ
a,(:J,eCA30,&@]-RcI<GE/a@1?b8J7<07Rf.Ue[fdRV2WG9dBb)8<>J4c/9K1^e
\(_XE@#-P7_#PXV;QS>B3,H+e(7[QGJY7HB.UbQOC&CHbJ#6L>=0^[b))^@3K9=f
L8&3CAJ<K_FUV@>6bZ2#3JKcH?DO]<4AO#68:fHJGd47&(])^b2-PWM7KI]V\W1L
EYdTf@/A6L_<X2/F,a33-L/JJ(bV,bZ@.F+J^N[Dd2(/L9Y6J@A(gLS+f/.K4F6:
&(PfHSMdR/X8PP#A_bX#.HXX<<D0R3DJdKL\HO+7HL)M[N(+X6@(Q@aWM7NE_MSE
:Hfaf(LWY1F91/POPb)PW?IIIbE7Ad&ADES1c-HUJ:.d9UE6fg[?N\A6F5F,^)F?
C9Xa2^VGSeU^f&eIEfIKH12U,GfZN5SPGbRYJL(=W\03JB2b1&8,FID_:HP:^<G9
5]YD-8,f0_XRb77);,aU-e(,72.bccSP;cSP0V7cQXCc+12KE/I@-gY:.NHc8WY-
ZMc8IUJTe+EL<d(4A.e->FFL_D]eG/Nf.ON-^0>=cSf)>+I<D0<O);SY9#OPU)V7
6\^C+MP@EW[Y/?4[f][Y=aNOCCAV@D8NO<7CR+@5ACS\]D&18O[9T28BJX+WK-HJ
9eY?a4=I2/CF>?T010=]c5IbLM_c6fEEf;P6/JgB@L-cK=T1W1F==1)\Aa]:Y8,1
V2VOZWZ(\cE4@]\(,K&9gLI>Wb6M^Z-KCKM_THBb<&d2[U?GKI@YdUSE]H-FVX<&
:adgRHcR_bZ9M@+HJ&Y4VXH,R7(gE:=W,X7e,S/bM0E^#[dSd0?d=fGSCV^FP-=e
IW^H@\Nc@II)]=</?2S_TA,P#(48L8cCH<FDD.K&BBQT-L;EWM/A@BB)E87RGRC,
LSY.XKG3:P0Z4U(;&T2CfZ9FQIK(#@M1+MDb2+^A.0+TARb/:GWRgJPPA7MYSE/O
.,^BW/7_FS8P(2Y<RT<[gI1L6g6C3\a<dH\N-13d3<aKgMZ01HO?c:#+BDWO^aTD
V;0\[UgaV>ZA@@L=M8K7fSM94VL)P/1+EEC(;,Ra><dDX&/PJb,:EN3)6D?Y9dQK
8g^@Y.QJ5Ob#_@OVQ]beWbETd@T+bPN82MWL_N?INPV9Q[/?_]5a&:<7g-7bV<[0
]bE9C?NKMF<47#\?9Z?V?;G]7,;F=f;d4R=LeI?a^B_.g,FQ40_>BJ/L7P>eEeb-
G<7_/d95ZMPId,P+V&fE2\&6&Ve)8M_G-7EgaMV:F#9gTcV4_:5=,00g_Fd-+\.,
LOOEL\JeCa2HOTAIA/WD-FJBZ(9Y[fL2,;.3VLY^8=FM1F3O._NK#Ff@6fUV/DMB
CP3WOV)CF0.@6P+0O,YS8F.0bLV<d^SS<5,01EW8EeP9M2KZ<FTWc\&N:Rf1OFUR
XBY\=O.a1c;9dTDK.#X/V]c+daefJGBP^G?,BY3Z45TUH(KT3Qb1TGf]U,E1?Se1
.#TM.-a/<TdC2(K3;A<f(MCL+gYRK;>OM?+[cV+8B9RgM;5QNBNg[.?6d>RL+5=<
>N9Pg@fU==62CT;4(6.M9B-T6M[e5;cB=R(<,=<3F7<;Z&,CSGNV-3E0efab,9B]
P/FJIER\TB11GXW])M1)(EJeC5.a+V_2g<.-=(#?AdbZF9)Y2#^\OW)R_Q#</bZL
:-ABgV+&A<&?IJQV8XDXR&POTBJG48-@da-A8#+AOAX7F9WBM+VKH,Yc63SeB6IT
e@I-1KDAUSXEKH^)TKXKMTa?#\YQ3(X,PAN0d@HA+C2fDK5<3Y8+I=_(VRO\NEW&
4TD9&)IeR5U<;7-J^H4,K+S4OML<KO#.#@)4:U[g7+/638ZgW\dKVeOIOS-=LR;K
^e],9_?<VV2cQFP/CZ9^0:FaBLZ4dbZ^?9#2]O+e8T8,G_?a[eTa]b;C;F6ZDLP?
80b+GF&2F0O]b7ab[d_>#:KgO[5RV?;2f]e#5;da=<a>.-T9bOJK7fO&#?bC@+B:
CMFL+^6QcIa;F1>F8(>8fV@cf._@H^[HC0N;?(UF:CE=?d@VUFJ<#.T_P[[C@45f
X[ca\O/,)g9&_=_SCT.5@@4Ef4R[dV[>3MGP,/IXWe6PL+HB8LGbH]53Z+=P_d&B
\^3/&05_+2Y.6NZ3J9F=4f-H3@0^bWg)Y(]1PLC^c5;RLf6@.;BfA+N=:_5-E:(L
H[-8GUE_?LWT6LK&/H>5c>IM;O4OL3-3a5<a/DB<ER.:6+UG8;6Hd\5\Y&.8BB96
KR0]QJH#7-RIJAQAP9:UN<XL-E5+AE1SA[e6X:[-1d_(A@;=44NF.TZS=Ob_Tb,d
.?cF/];YaBU#N[?_I9aFE@UNYOY8TENS8:;UePLe(\eQA5C:_K7;0MKCKf=5>aC=
eX6g9KdDI/?V5d+<.VHHIEEcd^KMfT>@88YS.A3-;731Q3AHM.><(8XH)^:G=H/0
S7fS&W#g5(Q-]D1Q_=.UYX)+XBL5f<6Ug@VA/A;@e)9QCDG0](;@21XQ@+PWCf-W
84OX^P^Bd?.A)-SWZE=QA5>d@\fED45BO6T#MeZJ>@#BR7Z)/0C):]K/@YI589f(
_J=Ke=9O64b2UcAR(.7)70O>E(N[cY#U2b7cJ/?>GVdc:?c<QK0Y89A4GT2E>DEX
EJ.A))4BX:5@:BL-8FYgdLU?E?G=BbY,BU@c^#dCg<S[ZQ7-+/QV>g\&ZJ-f=ZWc
Y5C^1:+^=Ke&9/\/Q_RWK63WX[R3F][,/FD;.VWB:,&.7C5O1EH\Y\EB#A+U,aT<
4&e0VDZa65)=^KJf2^0B01/<7M\L6C\X=(FUdW&MW@)SRK3C<M4GK](3O.93_]9f
S5+=8&CLI<P=b,,Re(OQ0A(5+cc6N6Q=H\T8@0VYNUObLZN1ZOee)X?^MZU=efBJ
1gHHSgL?4d;\XTVL.:A>;#[c7#;&5gZ-<MP(Y@21E(ZGJT^7@JEJYRJ@VGbU-dGG
/?G]0X<W244<:)PX:eZU;F^U:Ife:)FD(R4KJLEW<[aM#1aT#4\I)QSdD]GfK+8]
-f-/^+M#+eO[EC6AKGC5+(BSfZ&R4^O-W^WB[B5PV3E,))C#ZHS7&W1\Q<?.3(c+
+EgY<IB,2O34/G/gdC:5\VA@&99eO7Zc_Y5D=E>GGKQ4Ig6HDeEb@M7:,BI-&)YU
5WC&Q#K81TLNO;(FS,<4F/Ib,b&,>5MX6&QTa8P&EE+D(1N71ZYSRIPC^Yg-=9.=
K^44;0;GOTY29DO]A-Jf8fJ<\9<XFGVZ(R^fZV_:6d0]R7I^..(PH6,K5[.g&ZJX
Z<8RS)Jd__c]U,J_2>0S^\>JEII@6QTH4GOW0HPH([(8Ta(+9::OYNX,Y@cY.[LS
I:7T<\Lb1X34FeGbQaCdJ?dZ0UK:@_5gcHK(\>DC.<@#@1Z3EYF2X>SD9]ER7QP:
Y/dYQK(7IJ:K;38<9(-6^>.1AIeR-G@>N4].8QGOT8>NMGZ/dTXO6B-#?F179_36
GG3RP)>5R^@a=g@+&d3GXe+F_4CCMV.)=-UI/7H9;\4g.QG/E@0bT/c0b#I<_Hf[
DG;d.da#=+&#E9b/XB@[1M.G15X\>SYdeA_Ua^/-e/8/EILV-@3FbCHN=4@5[7Jb
cb<Mca3S_L\HFf0+BJFAQ<XOS/R<TY6I@Q=P\Hc7a@TM<NX^A6&S+/[[AM92d7R]
Y)G?TI#Q]WSX9_c9YOWBC@gX)\1>4GbWEcPfd?4L&:?4>A8K0L0?\OPg&7L4IKH[
TXc8EdAe6c+XVMS4D6HgRM.A^H;BD[XQ-gMdOR5F,:4@W47CKfY5#07S)&WBH;RO
.)4QO3E,2b/H48#6.QdAL-fI166Q,F)MC<_>ONHM/,4&E9_5g5H\eN0@fb7=E[=>
g+49I=9IRZMVPW<\\3C#T1<09XNR\5R-NfbH4&BWJ^e0SdeOMbMH=N3Tc5E<XAJV
(45<\KDTfcO0I67<B(R(R1(NJ0<SD>=MC#X1e0<-->E5FdNM15O+FX5H6bNLIJ,+
_FD4W.<Heg=X[FBfCGMSREbC++JPd7NVfT>5-@:L2SB32Rc[0#D;Q2G9XN-R9Ke?
R]<H1TMG.LffZ^6KC_LFV69JcID@=S9LZ\cC@JG>@V[TOEW-+MYTY0\fWCOB5U;P
YB7RZ(:g\<7d(JFLFM/?7\?QXe&:+?S+e(41(?fg56ZfW4,KKd:fB6EK92KRf<YR
=1d5>]+[B;]<Jcc=b6f9NZ)eP)a<@e<3J7UPgO1I_Kf--;]1A+aMfKNc0U3I3eF3
^Q,g0g2bP,fNVZ\1#A^5:37Z@P?>JTS&G5M^Ncd:J\Q^d/M^\g[8?PLafdZ#aU-Q
WEgbI2IfMLHNabS9XeGaGJQMSJ):g_A+(K6E46SA:=/EfT/Q38,D7D#<+>/e1N.9
-7\eR7[.7^15[M-2YRa3W>dT#B6Wf4f^,N\ZX6Ie+N/_GQ#,5e<c?R:O>?UY#f0^
[aT<aG<SNV/U.3S4JT-ce]QF65NL)V.T7EB<4QNQ#1T(dY9[bS\Uc^a\D1Bgb:UC
OZ5M9Q=7@?e.#TCeG)/dYHUc/Z_QMGb._Pd)KGH0J/_F8OWXGS\WY9-_>=Ld-:+g
3UdX,@\B4d2U)eKA\3KZZW(K2_e-cFDd:PISc@.QEI(R1(,XX0CWS80)JO290PU<
N:G^.JEe/e&cV)D+T=Dc9UdXS=(7B5<NH2IPZ09a1;7/e[XE>UEaF))O.]AST+FT
ZPB1TW)d79cP9)SgR3(c12Wa5&CL);\FDYS<:KB1BFAcG4NbL5?9:dJ7#4^Q0dJ9
U>HJE7C7f(gb0+,UJ>_7V2PDd?b5\FcWP8f5A3XZAA@9Q1RQC/C9ZN(3?NDcAD47
WECae[X3VYCVUaIQb1bAL=O/B@]2,:QA7-@B0KAYgNaaaINXW4TD6:B)R:LOI_]]
@;I]Adb3d<9W+G?+CKYd6,S1.,=L<VdFA)E3egAfgF/cJR(^SA;YdGQ\=PecR=A,
TReL_bQV,c5e(]&W4^2fHY::0\,f<2Oda132WQ(Ta0?8_K>YGbC(Q3HdU/UK\bB3
DXbV\&REaUeb,0?9K:P/7Uefg,a68\U30FZNQY/KA7C[@&X4QF/X4\dbe7X][M@\
Af;.]Ld3Cb-,KA9eXYI;72#1feQ[\A<Y)(=fYH8SYgND[,)(2&W_.E&689D/W)&M
GRDg_17@K?6,K+(7ZR1R2HcPb-)3T-f#NB\QP(LB+POTY[=01Gb-aU5?]Z[YE+.2
Z#RcC0FIH,OB;de<;Peg&XF2C<FR5C-8(KDf>)^[8I9+89]NO;H7;E^Q_)&>6)fR
7B0J9V(Z3WOLB^>-CC,78;=C(OHZSN2DC0g@MLIf1B,e9@dE1^Tg?LOCDgS4]M8W
GY=<)3RbB1IHT9,YfMaZJ&+Gg_YDR[G=#(QaJBaL/eH(3/7S00C)O-YV_(^XE4He
3LDI8CTPI+)De,7F82)Og=L+5RF?IKX4=_4ZOBaX.&@LMEUY=84PGJ4YaGP4Of9>
/,1^.:ISYb=G.4-IbCX3,()0f4:?_5Q-]0,d^Dd:F9-U.+g,816TL1:8fe2fAG.L
:X_]f/0:a=CRF19F2T^&Z)>(#Q?2@@W+/C)G]?9dgKOUQB>gaLcP1dF\f4d[S[\A
?35NV9d2XP9f53VPgA)3-E93NU;_J+/4#+J3#(O3T]fJ@eP62)[&1JK51-W1L\48
QB.,)._MgQg.TFU^e^9X2H8I@YgGcWD<d8a<dN=WWg-V#L@.EBYH,DP]S/CAZ.g<
JgNHO6H7BE=gTTHML4V5^<0OQ_L(^P2OOD@:f1^W0/Q3L=QS;B(2#F8Y)f7K<fH>
G_5Y[AUUUARH@S;a9]&Y-A5OXQ[A^aZJBGbU(aWFN]G+XTeLIcJ?98T<B4c0I,4+
\eNUM_;eUYca188fEgP8=b[#=dBc8EZK^R79e]&)L^QI]B@[/COF#GA0dY<>MR:@
(#3/DfXH@&>c<VCSX8UC(2;CP.[<)((JI\8^3SK/#]39)+O;K0IKP9EcAX;6\5/&
?2[.^_2;^GM5K&a(Y1de-I,=2CS=2:;G_=8[78GJ&INMe66^E4OS>Yc<QT^S)GM7
SWGPW]Y)Z#J>0D)gf8I(NY4Q<\0CLa7W_LH_L6\WGMOR3047d135a@3=\[Xed]YC
39\Cb1=,;gZD3;R)<=JCKS6V-47e+YPLA^U]R#4eIJ90]J^+87e(T#G3SV^d:C6P
QY#cb4JB]Tgag89f;&RT4@@K<=\\f7EWE(E:3=\)FPaCA(g37IMT^O-F7PSTB.5R
GAAgHgVRcS^J5[RC/S??(X,-KgBY<RdCE&6>N18?/>@fb)O)J6[03FbT52c(WM?E
EAE@f5f0OAZdeP+CVPT9B^6/_=^>]]b4d\Z^9=;a]4ES+3>4+>JTa3Icd:T[SRU_
S73W)(aK6bdUTNJ-BOD0Y[L-HUb;JNL7CIX/J_>^-Y8)1,&I[25N-d.gBI-3&IQg
g3-g8CWI)g[1)3JN:[H-&(7QZS;Q9J^<FOB-^e/e<K8T(B_.0-V[;6:]Z>/=U/2R
W5e<g0?Z:b&c.DK&:EUZ_3MQO(UX6GG,_-.&Z-?Q)g)5ecK#QfC[6?f4CfXg@=T\
@[H;N9F([6@d1?L<+QC-_:?^fUR0BH\HVSI7^^J7Y0fW95KC\Q3+.D9ME(A=_Fg9
YB31EfGG0=:\8K3HA:d^TVBB&<@6,A?gFJLB1/AY-ACY#0\J/DUf]e2\)TL)[Z(I
)Jg.:b>=9)P\C8EY&I0(5&_[SXV-gT/^Le:-Z8c884,PW29?+V+4X/HUfCBc:HeQ
#A5.5/_552_f0:M7/T8HN]EgM4a?eLB:\(&D(F?PQQA/7,GN=e(WG22>9,Z8\gcU
HZEDMgcWSD9WX(1U#YRRIKA-69DfV>eLW>d9eT<&<692]OF8RXFT:LW(.6&I2G.0
)M;?Gg<VE1U5U+bRA^JC)PEeG-2/&U@;XfB1LB7&1eeCa&daX+700-\2G_1+>\Af
S_34<B_FP;XMeSd]f0=61<4:Q+B4_H.E.HUF7^VSS^da])#HG?Y_c.ac_BIB+<E0
(+F=N<<4R&0D@JQAOcO>S>6K<]?g]X8]a:8G.DX[=-+KQ,:;-D<dU107@GYd^6:\
6I3[AB<;2FZFa2JAcLSP7Yf#b-;2U7=ae-Gd&Y58<JD1?E91FGL>f<4Hbf+2d>4H
fVFNE]&B0(,13\K\5@F;Zg0&_)fQL\G^8M=OgYcX?;_PY:\LGEJOZFL[AP,28&H^
],:(FXF=5ILXce^W@/DW7DM4.?@7A6>f+WR9Z(4C,]PN=<T66G.#Q>2)^Xd&+dH0
G3?MJc;8]_RQ+&QF6NVFLGRN&>,PO([Z.N+L3gXP=_U<&T4L59Y3Af@fL34\EL?)
>)DJ\QPET>#/_Ve8d>06ORB.Hc>SKFfG.X;ZHcEKY]@H0=/UOd;UX:2:6T-&53+:
9YLQ,H4-I=I1@ZP2WV5MWPCE&009DX7C-F6#K<TRPX;AfN__Q-?=)Z-=E9<87Q1)
?f@LL>_.\-]b?N>:aE+OM[UD)I=0\S>aCT_:-&fMMW5REgRY^#UQBL\WHC.0VXJd
/K]3EF]\W@DP(PZDgI]e,6H_[gNOZR+(QS.ZL?b,#_6;,(eg.W[-.4^5)7<IMW,Q
4I#87VL-J3fbG0bTeW0NZdP:=g_V3_M1OE5WbecMNMYg>]QT@=;S::L2]Jb&(IFa
8,O&KHSDdO>7K,egFd7-cFR>6F0MCO.f7NMSA]>a21D=^Y.];&We5@Y-S9Vc:?2B
2FF0P#1NL#_bOM0CQO;15VgR-5RZ0?c(D^N[H:cGa\g=\OJcf8<-M7Q.S/IQ:TE;
F5(a),f17OggH++^eQQb9fR+&+CcS]H;LBF&J,]T]d:Hf/1MUSK6BU2SIFS+,ERa
#E<HW2XT+(C1g,-5VQP5.>e8&e?3b;+W[fJ=O?@RJd?0HCE79:_1b<dd).QaI,@B
M-EcLV=YIN7[ebIeaTER&0LI#>-C2ee-d:a+0\&Ea>We5VAEIf199<)=M73W5+,&
f;Z@>AZ&a]R[G4DCHE9B1H2W-L4?+\=SS?>DQ4LPPZH?,,-A7Z+8&@/6E\NL3M#@
e;B.U?FPLf]ZIO[#3A:eXL><;fF<5#5)?YM+CK-f\>e[BOO+bS1&7aDP^:^O846f
:cS/19Z^KPC4FX/[a]>SF&\fNU6+G2+@:K15)[c@f./DCW8#P2XAPZ&W6I_Wg3fD
/b>+d#Mb;d&Z]RcX/];NCgP4JX0P>&ae726c:fVBN4@&dA1V.NeOOC3L2SB@Y64N
7QQ<4&TDY853J?U[TSZERBV:6:9:\;T]JPcOQKJU5R-]&+Z70>d)b5=AHd-U/>&/
=WI#F[E;Q6B@;254\N8e,E1cI[:^U4?geXb(c>B2;072+4H(Q6]a9DWLege9Z-4,
C@ZGa4,RO/)a-T,X#,@/Y3NQ6b1][#?PH[0=+[Nf,&YOQ)0X+VJ\^<R^_0d1=9<I
IET967_ZT90SNKe8]:8&@c;V9#L@7,Bc:;C\]e2HXWLT8N/T>#bd0KeHQPFJ8SXK
)7V+S\=).(YfX:?DFD_]QOEBfYY<06KCMD:8]X65^SQYV55bF[=5@THcV>R:K/)e
FVFUf]1cZ[K2g5,5aZ^M\OO<=4X\50=MD^#V.ETQa8^XX#dC9H]M[7aZXL++YU?Q
129,HG\V(YNS_dE;&bTEGc;bOMDE^E#R()eIcdXH6?[E+KW&\7CMG0X6HRaK]M;S
+dg3S[Sg_Q5^BI/IKb3SNbP^?U<O4CW15XCRb[QPA30f:Yc6\#0Pfa\H>H&d][0,
>f,,ADe=\\3D6:+cMH9A5<:Yf_G5^MOC;LScQd:a5^KW?OU^Q)EBU84+O@ff?Z#R
;W/G.2#:A,dG>4+g-S[B+&eCJ[^,[X7F=I6IG-HcAWVe8-:=&Z8:C3H3_)Y@L8O1
2b>@YbT,XK0ZC2^3-CgKL5bfIB/Qb5/HM6a\8J#4A[g)d<E5&+?CDBb]?C3JIDC\
CBH9.a)GS[F8:e6()LPW5^e@8@.=R]^8KOa>6&)bT@&SaKG&MM)X,BXB60OBSJgB
ab-^^5VMd#U4(g66?@=gg^:WF\#g,fN-b/48X,??O)_]eg:L2N4T7PT@5Y__)I#W
FB8Uc#Wcb,X^1]>BKd:3:=#JcC&-+.#QX)Qeg8DN+4M^XJDUSXeLee/#9;RAQ7I\
741S]F@U)V0_C).\.fE(cU(>4XO6P<_a<Jb4)XRZeH]5JgPFH\RWb\YVU,2YbMB2
C,_JaT:BT@A@5D4/:(UW<c1UK5&VRY@3063;bP-G>;D)Ne0[3QM]5PgWJJ3=g+>(
=N+94cCR;=8I@1_4Z8g-4&A_,M.);BSO,&^]O&UU5LG=F@\35Xg4]79BBU\B/JPM
\H:3(.MgD@-(?9N]PVd\GHII&Z&39A9NcG^0].=37bG?8@XKFZW8XDcWGB:8XDea
aY7ZaR>.]?DXCE2DWP<QYfcD=e=ABNLZ7:+J^c)W+JW1C6dXa;WPQ8RbNHW:6-=_
7.-N6)^</Z56^M0F:VM5+QS9eMBdE)>-554H[>3;:dBI;Iba]5(:cZ1Oc_[HH\MD
2f1Z.X1T5dc#BR<_)0dK&L_+3I)^B1f^6c2?+K-+Dc[?),PX<VJ3F40@fH;M?G_1
7J3R=3bLLGIfOV#>9Y9MZc[T+/]J9d9N+Z<G9-Td.2PH=N<,EO=S_IWEAebJ4T\1
P<Y[A;WTC]>[9I78.[.d<]F=WLMV[9#M7RLXEcC/1C(4>NW:GD6-fg>:[&Z)1.A2
HB+cW=@/JJ.4a4LYK];CU>eU/\4G#8N4CF30e[a:3^\A0#<5af\>WWFEfg.<XZ+0
7]VC)NeV1<ae[O?X[eIcF<^G^-aXaQT9UVYLX:35bK;NP<U)YV05JeBW\:RYO:OP
:Bga,6+B4E[N32?_4;?<5Z9Z=GBdP.Y2PJ+<M+B)0+3S]N;a&0\bRMKJgI(C^N,#
12I9<e15:f=W\JgUR<b,7c/e..^&K2N8#G)>)\?^ALc0].&1+HHF/Z7RWb3#@H@X
JK)cF+L4U:\KcGXVMI(5-JVP_88;#BUG^IS5\KH3A[5.aB#AbJ7dG64B\VV^?_;B
F:[0^07WVJR[S@<&DY^0\d8OaE(dA>LbX:#([768?DZ./KT17][(:;>gZ\Cf/QQF
&C;9>HJ-VOG;PZ5T(/b9S(KIAOX77f3.XE+U+gE\L,=Q?FfXQA<8c/^Ye(X&:]9,
fE:K6RaD_\W(.L.@ZKQY13N_UFAV0^9X;GLZe_[QSBgcOZA3].5&ND:Vd]H-,9K#
T]^5G8]R+f8<>L.+YTeW+F;Sd_NV#^[Ce9D:?0?>E6=92DBTOKCQ#J<6<e8\0YJD
RID-R+5<bJ^GLS\JWO)1SS[A4#>[0-JT_HJ4A[f+ZUCTGeWggZ(\Q2\E?CRE3F&#
<cgdCT0E_W/5R.AcKP1ROBCa2&@W\+eaRc6_#9<8[b6YQ1-#3;(8ICg58G@Z[DL=
+fVVN966:.28GI&e[HQW,GKG8fREGP=CE+,Iga>c#HI3D9Cg=US:0^9N^;]AP?(e
4VE[PbM)F\?;YP0X)3(RaILP,^0-3XF7@@T6?LORf#g.f[VQgVbG4QSS7JY/_0J9
\3g_EBV.d5KJX::XFYV+0;/XB\V-3gbg^8gS1^0VOf(<#6[W2201aRM7\5P:]fa#
9eYJT)&C-R>-=W#IPR>=g;CTdJV4F.N2=AB..[EIH?aZg?\=g@E]H0F9FJ_?fORG
;R=a<=W+KMgHX-WA,+7@NAXRFNVU?(Z&/JbAT=0)6BK>X3IX-:_L\_X/1<<2=ZSY
VVM0>XO#LTPRV?=JYH4NA8(H.7L6;TcKOU;FaP95[S<D<cQB;ZL8T/6aSY@]WJ6c
<J_I&.c)GH=>Gb#H,EB2dX^Q>96[(P(1,dGDNG]L_N(^T+TQDNZMK4E>^[KS#Q\a
&SQ/4A@PQL0Lb,+C06<<9KFQE09<T.P5W,Y))ZTY,NRbL)gBB83N;Q.R?0LdGcc5
1_bOOgYec,)1N(69B3NE7HR@;WURC9JdWQ(8_T5?YM1>5P_)QSVDHEKDZ2)^6V47
XW9IBZ:]#Z^DM<UN=)\&>3I5]D@d+RQ7Mb?AGHRT2_f_<b#Zd/QT.4P_aX>2UD/L
V(f.X&)V(g#_I-\LI=4^2aUWV??6d?(,#DP7_[IaUdL]0=,\RRP])Nd_@Qd<\5N:
/6OSeCQ5dXAO[QB)K^,J)9G+/dMR(U[)2TS12_?4.<2G0e9)#D^SF9WU^QPCB_:C
6UI[H\NXE(MRbAad4TWKb(U)\#K6(C2SRK#Q1?/BBf,8<7/=\<^<FUX#DV;+&F+\
[Y1c]WUOYP,@9M.N52PL)a(-+,1_>T<TaMdbP6R_IM>Y,,?94a:(0CECaGGfXfT@
af7c1bb=B,43KIbeQ]TA_@FUAe8^Se4:&(fU,PdN/gbAKag:.AE4gQ75Vc:7\(@Y
Y+W@#NA)4c42](8B11JX<OFSR4\4d>A05ebFBcbPOXU,QE/XJdHBHF]P]g7RYQ29
Q=O;W)\dN^O<L[;S\@I743LcT)fG2bE/&Zg1dC)#9FHFCb>Zed]0cIHB^3GIePP4
geB4LMU)]RP,K\S?c/Aa>AM]2W=DJbJC6+X7PJcRQQ2.Be+7\I@-]J4-\BZ4^U&g
4d_#437:XD+-CaD(GdPV>N;d8EKYB[>4ME1(B;1/HJ34#O,0\^>F&5ZLaJ[/#dDe
aDe_4VX60AI6PHOQFg,(0=KVCM[S>g7H<+2D9B+Z](AXSQ_3W>.\a[U]\\UNZX?d
MO(a@fDgMd&;K#5MTQ(5#N:J4^M6b)P=Tg41F+f5QbUVKX^0MLFeR_EHS)ZcDMU<
F>J><C?-O_=>MM,&8/R&/Pcc58a2YDB,)2]OIRIBKHB=K;8f]0gKIOF[=_=R]ZP9
&.R,N;fHYKZL80g6U2UO:2Hba;[MOZ_+T=;F<(gF0DS?-&/(Mb\ERK\(g)>L(@(1
CLNbaR1^]3_-C44YMMTVLX49A?+gg\BG/FHW/L&+GAaZ,ZL-MH7=a7)IY,_c?LbB
T5QR>,FRCQFb#O\DI/eXNHMc=,PLD&VNO9_gW-:><]5d;.<Ded0NT7ZCM[808,53
G,22-EHG+K#F2b8/OTa[Q4R<G2Zc.@).HOYfVRf@]MMAD<?--7R]f3Ie<@2B.gZK
]6YI.0]B5JLH4LV@DW5Nf+I_)]eJgAAF.BA8]?,OG84,W4f>.e3d2F8f.=ZgCZM5
Z8QUaH4OKN62<;Hd/9#CEGB,.:&RLQH;LI5[+0fX#7[NN8d+#g4\\AO?d11#E)NG
8KC7_FHK+FZ1,?<ecYQ0bfE-1O,A,<ZT3),-FVC8[9T=Mb:WYW73K<WZ;5SW<;9+
0=2-f-U,LMC[UF4_^DZN(C/OQX:(/=d.)_:8L?C==DGF+9?6S=1-g(PP4(\=Uc9U
B@+O#)643UBA<KNK2/Y?PS,ZT@e]@E)B,QCc#N5_#8BRNO;?\^70&We+KBCDIf,J
R;M)2eed3f7_>)4;C.D]5U668+8G:]U0>b]37)Me=c8f8((RGLS#UFc2BPJd/94F
C:XP@T3d@B&DQI<d3IdT-;@[N;cK4:8MeH?5S;<IQB-Z)\/]Id[gYO+79[?MS/04
OA])?_16_]>T3O;e)g[5@<K,>+;]QLfMfXA3?MT+-U.LO>g]bBS4UW,G#E:b#;N[
H]U#5^ESOV;2;)<6V,+@97R7AHYB#5Ke#?9(Q7C;4fM:>GZ]1ITeD_G[N]6LKKM=
:)_9:AM963-LY]fXUc-?gJ[9G7d)+0S=/f7KSIa2=9P6<&&QRHeQgfIe/E6CW3V]
:c)gK;EOc=C;,(J@c]9WNA3/W],-XdFg(]U7<e.BI[Y6+&O)+U,EbZ5:]/W]g\8^
ZcDP;aQ@WN>^,96#Nc1V04d+,96g:>.41WD1JGHJW5S>aI/[g(WC4Wg2Dc\UaW>4
cI_NO16YXLW;\YVMY6?NB&GCdA3HD(d\UJG?64;/WN,=ZaDDTSHC&DQMXb^M&2W@
.BUMU0QdQ.U,T1OFDQETeKPSZYFMBS4-9K4M:HCdD#)/DET1N[X)?fZ2NaQORMAe
]2O/@39aMe@cTaa4TYA(WT_CM4Z9)S5+-8^Y6<O3S_5VgT/_2A^/:)IX5T)IU72Z
I.3F]R4cHLe]YeC+HXc);0H=c@f1;_:2Afe/RU7AK]G/@5-?9bH1LYPE:77,aWf/
Z38,L7b7e=OLX,S2_J-H<T^.PBW59fUVE@&(6>N&>M<>fJe.G21aZcAL^c;GL13O
92T&[_g@X1,N=\f.UB:5LE=CJ<[F&L.P-K#L0P6&8(&LLF4M/7afR#QcEe1cAKcf
:1VHSe&\<YZZ?#_IVR_cG)5:NGcXeDLUK?]&RZ]9OTSe]G<4bHA?1e-#E5B#52VT
H@6M1NgMO=e#;X^^6]V<.f1aXO.\PQMcV#)N=J.&V.GEc(d5)RdSQ2aV>780S;)1
/7dAJ1<?NT<cCW1E>HB:<SbVa([[+bR=?UZ=d./Dd<HHQS95X[L,)Bg=g/cJBD4R
AXJK/R.#WH?M(Sa9Ka/^[8298)<#H76OL^<5JQd-IOW\]V7MVF0K9];JfMFd,>YE
X/V6_H2c:T;-dQPFJag+9B:A9b6.KgPQ?OC7+3TEB_4/.25&5^;27>J=GO\+O6/=
aD-=4Z)L,2ce.0BLF?\Pe/&X##?:;:]O[=:IG7=_0RZ+OeMdS7?R&&8>_:GH-dX(
X:N7FRdQTQL>cN+fAON.Y72fA@BfT6b(F6[:]HSOd.VY[<,;eMC=L]9VcE1M-Q6K
<ESc-8D))9MS@#5FeScV+DN+R\dV8Q=)G];0c79KYD_5G4PN2)<4H4V@+F0:>KC3
_2E\SQML<)[.5X2@>T(f8OXPS;Va6WPd1[L37ea8g1H#DT_FTd],<R@e]Q)_49Ig
.;Ze\.8Y96SH_Q4e?_J_b5KACDGb#PF_/XCVCfJeXEf,\dI)O)87M3]BFOSLWA=D
2O8ZBO[WE2L=JO^9+/Q<3<cd?>g7\e\\.W_SR]2(66)Y7a0c\SWeYTBK\a\K?9@]
Pb+JRV3ONNRNU(,d&AH<5PKGd(8_f^2LEO&[<6.K6b+MK&0M.YGOOFH3M[-;.3:K
EUK?66WVUc5D<APETb<d3HdeRg-@g=O@V)Q&fCKBfc1LcND+C9Z:V2>9b=18aKI<
LdCS@a12@3ccb7efQNEZf\_E/->AKfLQ;]/&Yf>Sc3NHDWE(X=fR25E,NZXJO1EL
P:>ANQH)FW\M@L(C<\\\Y@@_2E5=#aY:=:?+99e);>5AeQ.g\Q)=3aZ9[dG\/NMH
O1(-&+H,fEAa?U4:=H5I8L@PO-)3;B^^#PMO>+7[f1HU]M4+CL)P0B]K-J;SSdO:
(T-0RHEd4<P6OMI&6eaRWF,GGbK6_M+JHZ>&TRZ248D</2L.\,TZVb+18?>K+g-P
2H<-O;BKPSQ7->1cJ:JfYW\Gf?BKgde5S1aa3BDXCY+cPe??T^>SSDRGI_<4GLB0
S3P7#IM\6eVCO22P351G[EW(,8.4,>TU0O0Z3,ePbJ1?<,Ff-;+N-6135@98a@fG
IAQ=-B3=R&Q]aZ;<+Y.9MdHU0C-e#H9YU^.BLFaV<ddNT6?[I5TSS\YLb3AM75Cd
+:<7FC2Wb9fTFI,,:&(3JU#5XIF#OB[-JF5-6OE)WVS4URR;IJ00A/PZNSfXC3ga
79bPU21N1A)MINAegg1aP7EeI#&ZRPCL0YN#5>3(VC^JD7]7:e)Q@\VV#.g(+D(J
e\4ZZeD7VD(:CaYb+X]M8Y?B?41Y]MBC)#0HF8bO9PW-I\)2>U6e7@f#V/QUTV/+
IU=IO)9c93;d:L^RD7>6>GF,@S5YAc[<edag?I\[]RMbDU-U9f4@4b3&N220c++6
gc9:E#07=e@4[1bLD1I/K4&LZ2C2=A5:+#8fK0\I_#=I=K?@M;X^5>d>[bT5a-70
\T=\EMH62?XbW/4AZAM+BUfIX@=I=L.1Q<I;9FHWDS_8#G3@6=)58T>@3d]&MCY?
=Z#99?50b,D\[gJ6MC.0SOJda#A1+0#L,])W_UY>,Kg\MY^e5KW7DV:M<7DV(?g^
?2R77F2\4BNJQKHU-HFRF,O=\B)_VBN/]-)R\>QMcAXHbNNO/URgggZNG/RB]f#P
X;2,g0/O6,EN<5bKTRA4@PJDYBd+&FN[0)2MYf9REe33CfdL+T\9ZQKP_^JOd7Zb
CBDQdU^_fPD;bB5=)WZb66M-AZ7^[S#B(N4dD2>bI_4U^cd<;W?7UT:EMO@cI<dc
)M4Md>f?D/_.E6(GE+gRF,(AJVR33F@_AaNHC1-)fY]&@c#Z>9bH^&C(@Aa59W;[
S>T:4bTe^cH#P86c#V7Y3/U?.YATe;XL)4f8-DANeb&Z]/IL+@H5<;N7K[FC=\=,
DbKCZ/:1.JOG7#cdH7-D5H<O@O-f?XgJCf_NC4/:FI_74V1CZNbJ_W,_,YMf8^GK
<SIbS?I[GgY):N=AA\6\#?QAbg@^?e[Ya]7\5;LT:VSL67_9=4=5:7GZ7D1#8\P#
L1[VCK_FI=F=YW54[aOCE7LO3g>1C,_-U;_;W4^B3N8CU^&Q[#>fS:RTRXHcS6+6
F7._5X:JRTE2?a-Qa?gMB4C#FFSd@+VIg_X/8d)HWO4d3)S;b<YLCa^XN8_(JU]Z
KB,WX8Cf-Ie>_/U\N_++=MINA+]0-Zf@6QOGY=[PV_GT/#5H]G4C9c<.E]^R_41H
KVK,;949FfOb<-eTBVC<>QDH-TSL(4HccPCKeXCB=[f>L>NJ88T#43KEOI)bX\Uf
3K^HZ;,MXW_VJUJ:^:JJN0d/ZKL08KCJ<-#:+D#fO#FM/YfL]d&/Q4F4[e489<fO
4+=QK/KEPEC2N[P#Z_UgRUY9X97ZBPJ8=J^aBQ68N#24V?_Y1O3+4?&2b&KW/?=b
deaH67Z(H;LFe6M5g[Xf3FKH;c1SR,ZF,c04?W5(RNW.F&IG^#4(U(FM=G0d9Q29
aFT1_59=C-XD]]Cf[OU7-X?F:Z5<IgGIb./QPB4HA2ObDTc0\WS,b[1=HH>F+BD+
=J]F8b^>K1d<-Q]g=>fG=^XJBQ^F)S@d^.N(DKg:f6<H#[4a:f#LV#N3]ZbO/G=8
f^0>(<,V21A67.:K,E?f+Aaa]C16O<b3UZZ01SD&9XB.74RGId72:WG[e>Wb8XQ2
R\?KCQ#GBNS)-LNEF)bDLTG2B_J-WH>1L=9<T/6Q9K;G6UL_>a<F@MQR.MRcM,IZ
&9,>+C32G.\_08d<dC+?dgdIab)/(a2Rg9&dba#E+LJdTbZb&W>ed-_0LZFLB[0+
L>Rc1_POaRZP?.A1)Bd5@Ud7Z_0;EN9KcaMf7Y[GdCMUW?IL5b,YS>F/e))[a:ME
Q;6BGHf\UD2E0F+#+BD16+5N8+I>TPKTeJHZ-;(eEU3(33GeV#&>+c+gZ(.8IE7a
&2cWa6ER/1>Kb:H2A,[,W09@2e+)<b9JN_>D);#SK5/D^(5HE5FAA&XT13W@Q=)R
YffKaRg^gG.e+TCDJaA(RfdN9,GN&&PdcQX0])HCTa(:>9H-C@YL4[b#25CZQ/WZ
RQTaRD&1L,H2?IJ-P2K?JGCBE539\0e0DA:O?G918fUNMW8.TFC<R7>0VJ:_+cR(
U;IW8fT)P>^)>7bWc^E?C@J2J)AdBc,..^T](cNUO.SE@/-,d3Z&\34(9b<>DO)8
PC5^U=RZJ7./3LD&Da^F.K3?K>9P@I1c_DCI)TB6N].P-TURc=8<8_FB]bD[84<H
Gc[GTAS?>8(;@ZQ&0<ZE356D07\YVTE035=)KW<3KBZ)TWU36c1JL@.10Q<?C61G
FdA80Y1-+//HU7VZNUTGN=1;I0X()UVFD,KR1-<P<@OINV:5e^Y,E<OKMd.V@5Z/
@gJUVL^ONLfIGQ(d/\>@(-g_6F89D0O2:0&78]_JQefa#cI:1ZEB6GV&EYFDD5AS
@b]][d@F^94PD^L03I&g6g,Jfa]=-e#@,DJgL[9LZ8Q(.JP)ZTM9IB9+\=fNN;K&
87OM_Ne\,RZ2\U?bLBJJL]BYa=?>]AW;c,6DS&V-.TcdES(ZYDcVMKO1()5c7<VS
)dAPA[4)[&#QXXUP,_bg7W/;CdK+/,-NNP-N5XY]K>;[Q8<KZ@P_Sa4:b@&C\<2,
0U51]2Z2O)J0f:M1HD+<6:\^.S@WC(/\c)5T>#/@Ba&)aE&<:dfM+7DV6E[)W;Ve
3>)2TAO=c94GS)_[YBDX_3@8;a[(IQ.A]a[^76d(2K@6&J-b[7F#C3?JSK/\UWJS
gdJ_eD3cX,Cg=F9SZCCT^B65QTD=11FE,1\e];X[4GLP[]\X624\aYB-,HVE69VL
3>#7e<[4#]S1#\E1C[7.8CX)b;<PN6-,?+#@6a2_L,_QF>)-V.D6:+QX)4e/,M0K
O?BY>8?MXR)+:R9e4#GROe9[1:bEf<2,Gg&7?C[JbBO)._E,,O]_DU44X<OZ^40-
eT0<;ZLdb_NgWP(>WWgEK+W::QBAPFI,4BOPRICa]Fad2WeS\a,M#/G/X>OLf-CW
)cJF1+3]>a3).\O#>C4_\^/OUJ5J#LH5eIEH[f)G>bC3\<eM83]:UI6Y8YaCRM-K
4\2.8XHREI68X9Z=?<>I5>H<R;cYNF.c#R&[(4U^?cMJ>O&8L5B&eJJL_2=.2#1+
MZF],L8HV06d9M4^/DZVHF,G&V^CBG[S14HV[+,0\@<7ABKUb]KV3P[,d=8Nd7EL
E.^]>C)(&97^UU3PU<@0D7)R,Y+aFLAD,UVGUUIEL9@^)]:Xb&B>:1.D#--ISd@F
W+IM.bX#3(&M@^)I8,bT07b#OONE8UBB,5G;>>X]AA2Oe-,K6^Q+2QfX<(QM15Dd
EM8?Q):e&BVXbV#79MFI>HVLEM&a;Y(V--9/EM94N)L:R<Eb190:DK#=MIX/+3/,
,^/f1P[.35:R2?69]aHIH0YWEF4JG+\).Y;E+aX1VG9cG6.ZcB_J3HM[1OCD7AN5
4_>6aO009/H&BAYa+[EYLIR&D/]U=.f3FYN,aKSDMYJ?>4d\;SHe2OYe6KI[7B-A
Sd&U^3^BZ5VE&dZ9VIbYNY=Y^U3S.=V.6SGN^FYRP][a7<O]a49T.7<HaQ7ffW2E
U(Q-5Z,gBUUQO38Yfg<_M[JgD]dE5O8LY4=OIIVPI^MJD/<J+H13H6JBR0V-A^KB
1^MUG?.gNCRD:3E+.?XKI\e]XgQKI)GFJA[4_SB33;NRP)<R4<;6gM[Q>Kd.S-Q\
_.ESLC@CW[#\=N[^(<F,SQ<+35&D_YfC4CC:WI&;IV[:b_\Q2/&47>ET>2&=VLGR
]J8UYK62Z/7:FcL578+NCFYQ(1PNaOD<VRN+fUL#Z&5WLXR3X2c3;)9B68bFU:1a
X/Q@:Q;UW2T:#V[SGA@H0^#==1cdO[,E4L0+A(0Z9^A?G[NF\[7Y:O(Pb05N@XLT
6(-cXB4cKX8Lb7,EXKF3N9K^+L.7,,>Z;ST<?Pg(&6Df2G^2M3YI(/XY?CY.KCN<
\[ce:2g6QZg:=HN4B&7UW@]bZS&VD@D[FWLICT0GP.a.IL3X8L33b19TKO3:(a:(
#f=]>1\,W5]IH.456121)UfL\c:Kd?WH,6Cd+9>J,d_1DcL#L<MdMg\^g]?W#6e@
Wc#=,OSI\cK]O@9CfN6WK@ZROg)Wf21^:36Z?bQ_<(L8MV)_:X+<<aY><SY)QfF.
>R\S@OfKTP<SIO=+9,9+0A8LL)H;eEQ(&C8)gK73/>VA]_<W]a2T:HKN,fB_;Zg;
;2)[ZeDX^gC<,:/QL2c0,NH<9^d23+>:O_gM/&fe89WIcW_Z2TJ:.HYEO[/14<EM
#Q.J<CLb1MD>eB5;5d\S)e<gUI?DQ(NIMGK>P.a0^5gEP0J\bGMFT.CHcO6&g>#e
FJVOR03e9dI0R<_Z.G?#^U6X9gdSDKE@JS2\O=+NU32[JY9McHUKYLGVaMQMd;VX
P_9,IKBVDQPcN;_8-Q_+\JCD0-RUV93<0=C/-C.@M5E^R:4IH.S4:2WQb9(2A=0O
X4=\[ISV]](2=H^a51e5<X_<<_E::/C#d,,E+1#](+9fCaXE,BLRI_6TKFNbNR5,
C?bYT0T,?:4M->^f<(VH#LA66^IG;8UE89/T:c7SY^X2-.+AcV+KLCeC2LNCR1&:
a-BO_H@W?PQ^gDW;^3U/g2.b<VP8\#;2I3Q]YeV53^__9A&dEf&_<(S(NaO&Mb-X
M)RB+QaK_[+.[EN4C9S^1#>@(VB>5_<D+g4a.BgA9EVEeEK:T5GDH?]LLNA(BM8(
e\IEH&0Iaf24<W,,ZPZ7b_[aK6-V]AfEB8&GJcJ5Y@_NK2]Xe.;]QdagSg7O;\WK
5VU#\I[=.C^C9\=?1PQ&DT/>I3H-)5.U^eQ_:Lf3H)=<1E1Q<RB?#f6ILEa4VD/K
QOM-GK=bJ[D8XV-)e\J)7BE.[B4C@:_(ZN_df\c3e.fX7<:c8<-E#3J6P#dOCAG4
\eY^]K[[FBY?cI\eVDeG-UG-W@(D/)5QV_VI@55&/F5&>R=VaKdTXE&_g?J8C&<:
]VOZDTU]+DCHfM;3_2RaR]fCUJc[.;BKbTB?V6@DJGK@I-eI=F5=UFVXOGMSS-+O
S7I)Bd4eX6I-V07=X73L9SFeHQ0Zc?#f4:Y@WMT)E^@K2/<FQDId;O;4XCRQ^B;]
f0JZ:E-;G=F@#2R7(D5gVW2,CM9f^_[EbB+LXW8])UNTea91/9.PG#BfUBD8;A3d
f/Z^WWK8G[DZf3Fg_DA^3]Hf((d#-T+M)_/LOI4G@APTZLE]]fIIa+4@F>8?f]57
_L7\g+b=;^_<&HH2[ZV+X)EMN,.,T]fBIZY5FUNN]H:&ZI5YBWC2O;]e7;,Uf?KU
=QF85@\\gSKd^EG:7X\A2Y.INPH<@L^=gLD#X=UAF4Ma<bJ>YZR4KZ:6@[=SHN-;
1<8^??0C^,JT=Cf,f6TM\UCWS(0/13S<PRDeW2R4G42EL-^NF,PBT;=@?>^NQ#G?
WO=+;L]dbDL?F<FE/]?bDHOW2(]e,>ADF/\2T;JX1JDC06HO6LaQ.P_.G@+@D0Ka
6S:B[2B9->G?QE=HeEH:JJ]<CfVICIYBF=TM41CHB7:)V/1M:61X8&R92VE?[W8B
DT924#S?=AQcSFUAN3,;>T2;b^FT):^T,RMO>+0^)U,gIf7ON)#/RMagW2?^H-5N
S8_7,[3Yf#]/M29RC+ScRC@_;M7X@/bf?bbEb#.TC[A:B_5a6LE>&AIbTEY76Te@
D\.2g-7<K,QNK)XAFB>SOT^).b2COL?L3GbYD:Y^HfET^^gbYF/L@O-\(UX-@VUV
04-\]?&MM#;PJMD#DHb9Ig0.:MI1V^FSG:@g9:[eCGZ:2+L=6&a0K?-_B9(4IBMd
b0DdQVYAaR(c>Vae<^)-,SNYO9\YK#LF3F386X)X\&gN)8A@X;46]@NHTO=)VTP9
&dgJDFSCP#GU&HPR.YPTZVa^3Vdg;AMXdO5DRXP<D9dP..\e6\4/dUS0ZNC=49??
EY?7A2+G7Y9<VYHeWP=+;1@U;e2Y&f,bfA_ACTP+]SO2-,Q]GB&Qae>OQ:OUWe6)
TS7G/+SMc[0C5)#R6D_e+g&FCJ?1A_2WK4/,bECUcMR_487cMGQ_AJ,?KW3[LTA0
?OaU+TP?(PR]+c)dH<AG>HBR]+ZCJ6=Q:a24^e#)7Ac\_;-F?-S9-SO)Q&YLT&Me
)bQAb[LOXWSG</GA9P1Fe+Y:f:19(5VP6J_G=A56YXX4G,SB[0/=V:F\6_+V)3,?
[ZD5S4:]IH,JW/eG^_;GNR.#:P^<M4T@OJ7U-6YG^Yg38O775XEA=&ZfBUI5eC_2
)g9Y.#S1-9.+dFK#(.CgB0VEFJ3a_(dD?LPI,CNVZ#b?5?=YEVKCKc<PTe;[@_e=
V?;eH;QJV0Gc4LRcS)4RX:66L<FU#]3-C?>Ye^#&We5;e52.6MS:X+I?DZLf0J1K
c6^#@aN/1NS+G.@ZJg-:PQS?7a8;9gTPA;>4UK5ONVO4c.e8YL16&fB+TgI=^NKW
YAO?L#;>3?>&LG8Q.ZbYQG)9GNbb&)1M[/\-V2SN76g8(4ff,U?W(ZEFXV]Scb]D
g4aOAWcaHE;\@F)0O7XLB[JC=Ub,()bH0\WXN9?Nb,WMDOH19[/\8.c[&_F@d,W1
;eZ<+&+;J_e.@)f_egcEPCPP=-K)FW9)>#0dYf[[96GEVCE4;1eLLSTEbWbATJBD
ee6-b6ZXG10/5&E=]47)QZRFHd]-=:U-#S:NW?;)JBf&Me\:3=-]@?SEJ(0:@-<X
4-4[G0PYEa=JE(4a-KMOC^R:\^FDE<D@c0WS.;R5O:4[P0[(QPBACG/[VN6<+fL(
B6@5:7SV(XaX/@DB.7W[J/EZ#bc,,4\J19KT=W.1:&#30NYK9X(.Q+\6eQg69F]2
MN@FTTg8R.P7+KdRAO\Fb@9#caC)8d)HP#]/1-A2>]<5;AAR&#CO2&YSZ,;@GbE8
gSXd5O.7#ER=32DVB0.^d=N)C==17W7KY:9IH/=L0K^<Gb_G&NXA>H+E]U-DPMe^
c7^5>@:2HBQ8L?Xg/+K#P3[0=gV\Eg]L[=H6UJQPaX:?BNX;CSSV&d97,_0>Y7_X
P<R8@/N(g1CCbWIPO?@3D+&@Qd\:].f22>7292;&Y):FAKB,1-#TBQ,OHIYD<b0d
69+LQIAP?I,;GGE7Y.ZZd8cCJ&F#K&:Pa[_/?#4;(=Re#Ec4&IEaUgA&=c5>?8(<
84.>CX):+]f+?W+JP.Sc\#6g+Ab(aAHDa2#5fT\]2:9/L-5O>I?A#(g@,PQ@]:MX
923JX,^85HC<0:WD-f,?I,WGS7;GJ4R<8&c1dBQf<Ua6,eU7F:b=KKd:Rcc_#6QC
?78F8<A\a5X_bM1F:-2_9AAcCcX\_D5L8,<R5Vd/BK5^?f^UMK]-,2<T@/6.CO9;
f(e;DEce>[0ZE+2TfbWC;FcX2\EdVR,A]XTJBee)@a0:[8/]@I30,.AdPAM\dA=6
E/#VA)U62Z-7f/,W/\\;4bfHHN)eFJD[O-9EL<L03R7BQC_[ObC]:fJ\5RK=[?/f
K8HOR.9\FbI9P?XL&V3g4<6?-_G)PCQJJYEBFMCRL6A9Ac<>P.)/Kfe(<f<b(aQc
^?V1TO5,bO=Pgb1e2(\63O821?X3<]M,DSU+RXQ@3<8BEMR)c=MC?<JW@71XNfC[
D>_0P2HNK\:f;_<[8LWSMf,cFSI1Sde&Rf2QA=Q@OYACb_fEM&?;J_Z6>9B@^cUS
ML7U\:&Y)PL?,fK@5I3.OfSf(9?)->.6a)=Q71&YaZN,(FEcEI+778,[F6=QLT)J
8.\5F\+)e1O@/>?cJZ5PN3Be9SB32OOEN:X(H)K]#aY-F\Scg<V\+[)aK8KWd6:b
.(O1cNF-9K;JI21f[dYT()QZb1J,EM]#TYQPMCFELYe,6)ANa.D<d0I6QY0J<8,.
_U9TH6G__WA/>?-N9QP,f&?1BK8,7N]@JZ.JdVeIcHTFMb:Gc)g&T/(<ec#03VB>
XOgH#b]RAbQ>1WRDcO6c=c.EO0cQ=L-aJZ_G19ggET7@Y5CE9<e[O=&R7VJ+dM;Q
)ILcMYQ>^02GEF>ga.4/&3W&B7_OWI;0E5FJOLL[VN&:cJ9K#@)WJ<>X0g1]@XZT
@<,Z.98b@M[;5?(N//]Y/eI/?/ALeY5b<.YI?6>?-5;bJ:9b8Q&29]2f()HP=)MH
^#/3(;320D4UW.;R1VP<OGI@(5bcHV38Y3FBOO2N85<P[g4d;5@F.U>E)1eZ/ABP
UJ759[eZ[:4D<]_,,cWH;CC0cXd<(UQdA5VMgKIbD=;RK/U^32^/LU=9a3,E[-GR
J:0geWRdI\Cg0-EM+8EM?CLF/BB#K?)QIW7:GV:V<9D;9OVM1@cZFBKfVR-YE(Ba
9ab+<C)#9KJ\1Cfg-#7<Yb>?gC@+LZB]bHbac9W>8C,.-ed:Q0HgaffRd?BF2YYg
\^@\(MQ;BD[LUEZ\((,QT^9A+;&_4IX-<fY-Q^Tb9(TKGRQC#<R]0BYf_1bAYZDN
c6Q7CI2=6]1TNTSK^K/eZKL4.D<@Z5(FaN9b8W?B_[7SUb:AD+UfL,B)KM,\]:;e
R86Zb>;Ea4]d&DD6I2EF9:X04MKWF2PJ\,#B.;W<\QCOSdP--JC7^H),]H+>NK>Z
bgW)7-W^:Bf61NZ:bR:=2VR@SZZAb8._HLZIeXRI#R;;5^85c[:eUO7cO0bDYVe]
G)ZA(Y]QO-^<Z/JZ&GO9]H+M@fYKg6J7?5ULMQQca_PVJg\TSeTD;8VYU>P+)Z]J
F.-0K[Q?6I8K?WAb6.WOVD3U+WPYLWPN/?>Ff_bEOg\,1.c?aC88KCgd0f>E1TgW
6A3RZ)VBSTNUaaXf;SHgZO2.>ITSZU5PGA]X9VEJ_B?+\eHZK\UPQ=Q9EFA)eP[M
4/-4YL6f+3QfPG>E,?@]/Z8a)-9Z;#-O[J.BX.:_5M:\F7d-BZc<OdOf^E)gB.g)
-S8d2OaC,0L=JWJ?YCfQC8HSZ61JYP&8:TB1@adaR:=WbCJQO;H[RKI..0)8I:F7
,]1J<BNI.,EY8HIN?5&Bf9GZ,d(b^42?9?KRWUC2X..@U/g[-S4PG9)]Xg?;439M
NbB-ObB,\c-I-AH?NS^6OHF:#/UZ21>#1UMBg3BPZ9TRVb.>E2ZRW\W(WY+Wd;\B
&9R^A1,V2BYCAX6_5^I[EFRLBGOaSF>)#N/F]YPPU0P#R6c;L:gA(V6MS;ReaZ85
\2ENTSQ#Rg?3OBcPY)(5&)4ac&_[V_^A>ffP_;Y3-9_7M6N;cT^Q:6F5GU2Q]M8<
g=7QT607)2YaZ83IJT+#.NT[WV?-g:EN+MbX_9;+/;VBd8-H=.9cVbd7Ya.IZ9CL
Q#7Q?2P+3R<<JOF2eaL;U.7Z,>17@EaK+g[0Q=IXT-YUQHE3-:g6RRL8bP8,#[&^
_?->7\bQBS^-5YYV^1b8YPLV\Y^IJ)-CFG0-/Eb3e)#bW[R=+V1EY#6[?,V5(;4K
P/gfC+6]EO0;)gfHUD1TQa5.YB;7(O2E<_c1a_C6X+9A,8P5f4-S=X,41PQ@[0N#
fG;E,C:L@aE^@@@.OeHac>bC17V1H]<BGYV:4ggOIY30S0B\Y1d8g@QH@2>)219?
eW.S#SZVc:..R\O@I_U^44OBe+AP;L\F-^\99S3_b&1M5VNDa<]\I[UVDZ=(YZO2
^#dcS1E]E9DdWVKFP/]\(@(Z)LBfZaZKKL1ZOB,8B\Rd?MR:=P&:fGB?OQAH9;1.
X1LQM.A9:6A<Y@C_7J1VAI)Ld@R4)EKe?b(K:RDc5e?)8a&TT/dO+>3ONO^2]\Ya
<4S>cUGU)^Q<.L-edgVgR\Y=aNgaUC((FULM;(-[2P&)2/fJTN\5[H;]0W/g=S9Z
<;IZGQb(D_IHD338DU7B?JfRPSP@][0:;cJN<+[&bXTQL@-U^\1V#.I,AIebK?);
(A\W+V50,\<Y8&DI;+;1W\SA&U3e]+DRR6&F;KQBG0gb4f7P0TB5;FFFMUP0\UT/
,H:0C:A)2e0A8Y&cbR]3C2KRA6B/(e-/GYfU70J]FZA(&&&-b[8W4)KD5Y?(;PE&
72CGIF=,#39KdJD^&:b?A-IPYM,(5)&;FgNF@7O18TK#C#6@bT2/VQ7-\,fc0EE?
(Jaf\a[(@6^Sa,N;W_C5UG2R;LY6]D<(;VT+0])]Y:9Q=U/T&B?[0gPBAY@d::V:
;f1-/_:ER=G^B8bV+d:A=,b&6HWIA/7W_H#SC#?7M(..5E#?=4A.DUT8>=\OCgCF
^H7O[?KW0ABY=3,OV<^S9AgTU#W+W[HCg#GAYA50CY]=#XFENWT:3>C/bPZ[K5AA
F6CKg3]+[K)8CO[7&LIZfI5O^b)WU3P+]DeU>a?@<S)Y,I^.9HXF-c<dQ[>+@&LX
C)eJPaQK4P3N#QVF;MT1:&/3D3b-]:MU^?gAFJ2Mg=Z<A//(^NJQR<@0D>/c_36S
>>0XUB+_HM4\:?^NgceF;bFH/8&D:L-L@R^0^W8DX:@cC=bgY@5^/?7MeI7-Z)\8
]ca&???Y2SK:ZD6Hg_5WCZf_HY6NKT>XCf^R9T<U2[(=a1SA_/N/GIMJ+NZ\9b>?
TJJ9)&@>JbUgR.S>;NUQcTV&]8+\Db#I2Z6P.301>GT3MbPePZ<ZD\V_-^AHJ[_7
(V;G_Q#C2[-_Z&>K1^EI>/^]e9JRbTJ_[>MgN]45Z[F99fG)8XD/FW,CJ&N=E-(#
Cc_ORI3=[c\VY#X?-EK=g6DE8fc_aFdI,7FX86_?aU/-3#a?5R[]VC_QR.#M4TKJ
1?Hf@G8eH?Xc1]G-.UR=8_T4U>IW753f?f1[YeCda4?EA+e(OCaU5Q#8?U.SA-WP
UX\YJBaH;b<Q@R6IJ65aD_/1Z]:RD>0S7BS:6KMK5C&C3MP<Z9)JN<7S/.d6?PIR
0.X;RQ:;4RG<aB>>C3g7=IL)Nc_A49+\G[2Q<+Lc/+4fJTJ6KCdR,f-Y\&3F9_R5
9Z\ZY5>5_\2]]VB4+M2-4e:EGc2RYO1WEO4g3O?:<QC/VI3^,]F3Ya4\]<,:ggGS
6I0VE_G0@9fS/S,L5N5]TY1DN8RE.1B@@3^0bF4Ca>aVgY#VYZdF.;;;=e#93d-&
[P[<A@U3)RA4Oe5,C9FY8?,dB2aN8CF^J8E,dXQgIJb7=^(PTc?D;<^\TYHV6b94
+L>-NP92(]-E/O;MXaObDgRD1c;b[^E.?Ab/e,9_(D:\[LT@J76/W#BEgZ^VJe[:
X=):E\2(8>,9/,Qd=M<RKgJFfEYHE/(5[E-F(U/H]62KJE.]]a;PX2d:]J#ANO?R
c3N#;.>E4XRV[+7A8MOc;@PE2=6caRY&^b]+S8J]CVXg#RZ/J=0[>XTUNa84.5aI
\&=5K:4)@@aXBE/^/bY:g_/G\H>(Y);)/QbW]acY89G2..^=g1JAgd700If3GCDM
O8/-TeXTS3.K<e:OeOP)9/aH=I(8G=2WYC]\S)3CWT-?A6ab\=T@2aCI\EO-+-V7
][MV&#>[G>+6IbFU]\H]-<CEfc#<L/\e.#HF:f;;N2TA6S7H)Y)96-W:QEF9])4K
XR.ZbXaaQ/WHM03-A@VXY(^NC[135+A^)3RG<d^)IX&E-A/.e4Z5<QZ/B7MA0IP4
\@(-W4-O[Q&I69,e0>[XV>.Wc1MU/YOND?>>KF&;>6B5^ZK[1eWF)ZAT.&US^VMf
O1ARMAQ3(708eg0_4=,BJRE]#b928b^96B;/W>bb-:[]c@VR3a;?^_Ag\.J>5S>W
X-:W\RH=6b9a/\4IQ#(<IAD@_O;-BP6R7=bD]SS3]K<K8ZZ)9TX&TS?1DcaeIFPM
<gTfE/3I1;+b<.8#J,3e[:9Ac,gQSKA_K@I]WYNIR/SR^\DZf<d080,:HPH:6GO>
-?ZTeg36Bf.)_9a]\;X<Q#T0?:TaLCgYA(T>(a)c&&+(c.>-8\X3&.2aZAfU9,MZ
.:#^BcB.Be4P+1c7[\LYCF]VLUGDYLaTgPS?T56+?8ULe5#EXVY4210cKdWY_>NY
./<;Rd+_;;Ie3_)UI\acKAV64HVS0<KfCL/OZ7Y,(,_=#B&A@QZ6+T6[Z@K/F=D3
c-eI\Z7&JUF6(SO:@[S6W#H5;^YgIGY&NXSMBZg2(:fFcURQ#NcZL[CCV,P)c;6G
Ze4NfKI:dV76_SD3e1S(V-)WYH+Tf/4MOGMTB&7271AV/IaNP.H.V\\34+T&81_Y
CL:fXB\(Ege/5?+>_<3ZQf]6)BZ4V,[EfI0>g[b)9ZH?L;S]]3ce5(3b;N:SA>I+
7CgA0[=e0#9EeKX]R8N9#7=(U5U?]=PI7IA,(I(0Ne_4R6HF/586143bK3LU=G4d
573#K5J7EK]^B#(ga=J<-WCZW@7QE&bV(VE>(LZ64H6@\Xe[Q@-T7(c8b=^5YI\2
1A^<WK+0Y-YSKf_J7C_fI9KA1V?E#QcgO#U9)V0-KCVKQXb17X0SR\T>E/6YbBeS
KU5H-ccaM8UR:C0KM4W&FTY>O_1,5.V(Y512)S)Y0OBc#d+O>L1=fWGX;[G1WMKe
Ia6/\7DCF8EDg\?2?;]=BD^;]XPG4Mf+:9;<E1b0QA=()546==YV#)6eBI5F]9VR
234AC8Z3>E.Nf/&L;/9[Q3YQ#dX;]ICM,6O_26<7HDI,;F,>W:7a8?MIbX76/Z(W
E(Z_TYN1;P&,]/AD.]Ia>A@MB]\2CDZ#dG_@/:K_3c>Zeee#f0DCMW;9PU\L2:&K
E]aQLa/XO@+@;f.+_#J-D[7(UT=Ve5JLbK?J_.b5H(NZe:I5.\8HLA&T[E54XGBG
?RTIJ;MG.@//0?&6d@5KTZ&\9(S+&Z,M#FBPZM576,&gfN;=98Dg(TJU(I?VHB;a
9Q5M&02SVLRPa;gF[Q&=^3K-P;4EgN]>e;>Vb[a(F1^(4K#TbQ\N.L]\\:g?3DM[
XG8LD2\@G?\94:0a\PCAgVR[-fbc8>cReA]O39EG3dOfcNRQVB)2[c@[KLEb#&@7
<e_0.)/f3#]Y[U.__;#E0?CG6\6dP?_CXUALC,_CLc:FW;0OdYU]6O1Z&5?(A)@1
eJg7=cLQfZ;0?RY.EDF2(ST^_7F)Y,#I)TG\XTZDIM_B>DD/XS]80NdGg47KE4@Z
@1H>bUWe?[aYL6:5>90MVR&dfXVb5]P==(;47XO382MDaKP^7dY<;)NS<CL-G-=@
L&?R8;N^9G<VB@KKMC7MVB(FM]DcPG+M\XG(91.K9^9e;IW/.I<EX_1C0NeT1QX,
=]U0Y,R8+:/NE_EQ7Cf87E5aOIJ)a5P?JCZ0UcU,U<.AWaUd^YMgHV1CI$
`endprotected
endmodule


// for spec check
// $display("                    SPEC-4 FAIL                   ");
// $display("                    SPEC-5 FAIL                   ");
// $display("                    SPEC-6 FAIL                   ");
// $display("                    SPEC-7 FAIL                   ");
// $display("                    SPEC-8 FAIL                   ");
// for successful design
// $display("                  Congratulations!               ");
// $display("              execution cycles = %7d", total_latency);
// $display("              clock period = %4fns", CYCLE);
