NAMESCASESENSITIVE ON ;
MACRO CORNERC
    CLASS PAD ;
    FOREIGN CORNERC 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 235.600 BY 235.600 ;
    SYMMETRY x y r90 ;
    SITE iocore_c ;
    OBS
        LAYER metal1 ;
        RECT  0.000 0.000 235.600 234.760 ;
        LAYER metal2 ;
        RECT  0.000 0.000 235.600 234.760 ;
        LAYER metal3 ;
        RECT  0.000 0.000 235.600 234.760 ;
        LAYER metal4 ;
        RECT  0.000 0.000 235.600 234.760 ;
        LAYER metal5 ;
        RECT  0.000 0.000 235.600 234.760 ;
        LAYER metal6 ;
        RECT  0.000 0.000 235.600 234.760 ;
    END
END CORNERC

MACRO CORNERCD
    CLASS PAD ;
    FOREIGN CORNERCD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 235.600 BY 140.120 ;
    SYMMETRY x y r90 ;
    SITE iocore_d ;
    OBS
        LAYER metal1 ;
        RECT  0.000 0.000 235.600 139.280 ;
        LAYER metal2 ;
        RECT  0.000 0.000 235.600 139.280 ;
        LAYER metal3 ;
        RECT  0.000 0.000 235.600 139.280 ;
        LAYER metal4 ;
        RECT  0.000 0.000 235.600 139.280 ;
        LAYER metal5 ;
        RECT  0.000 0.000 235.600 139.280 ;
        LAYER metal6 ;
        RECT  0.000 0.000 235.600 139.280 ;
    END
END CORNERCD

MACRO CORNERD
    CLASS PAD ;
    FOREIGN CORNERD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 140.120 BY 140.120 ;
    SYMMETRY x y r90 ;
    SITE iocore_d ;
    OBS
        LAYER metal1 ;
        RECT  0.000 0.000 140.120 139.280 ;
        LAYER metal2 ;
        RECT  0.000 0.000 140.120 139.280 ;
        LAYER metal3 ;
        RECT  0.000 0.000 140.120 139.280 ;
        LAYER metal4 ;
        RECT  0.000 0.000 140.120 139.280 ;
        LAYER metal5 ;
        RECT  0.000 0.000 140.120 139.280 ;
        LAYER metal6 ;
        RECT  0.000 0.000 140.120 139.280 ;
    END
END CORNERD

MACRO EMPTY16C
    CLASS PAD SPACER ;
    FOREIGN EMPTY16C 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.920 BY 235.600 ;
    SYMMETRY x y r90 ;
    SITE iocore_c ;
    OBS
        LAYER metal1 ;
        RECT  0.000 0.000 9.920 234.760 ;
        LAYER metal2 ;
        RECT  0.000 0.000 9.920 234.760 ;
        LAYER metal3 ;
        RECT  0.000 0.000 9.920 234.760 ;
        LAYER metal4 ;
        RECT  0.000 0.000 9.920 234.760 ;
        LAYER metal5 ;
        RECT  0.000 0.000 9.920 234.760 ;
        LAYER metal6 ;
        RECT  0.000 0.000 9.920 234.760 ;
    END
END EMPTY16C

MACRO EMPTY16D
    CLASS PAD SPACER ;
    FOREIGN EMPTY16D 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.920 BY 140.120 ;
    SYMMETRY x y r90 ;
    SITE iocore_d ;
    OBS
        LAYER metal1 ;
        RECT  0.000 0.000 9.920 139.280 ;
        LAYER metal2 ;
        RECT  0.000 0.000 9.920 139.280 ;
        LAYER metal3 ;
        RECT  0.000 0.000 9.920 139.280 ;
        LAYER metal4 ;
        RECT  0.000 0.000 9.920 139.280 ;
        LAYER metal5 ;
        RECT  0.000 0.000 9.920 139.280 ;
        LAYER metal6 ;
        RECT  0.000 0.000 9.920 139.280 ;
    END
END EMPTY16D

MACRO EMPTY1C
    CLASS PAD SPACER ;
    FOREIGN EMPTY1C 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.620 BY 235.600 ;
    SYMMETRY x y r90 ;
    SITE iocore_c ;
    OBS
        LAYER metal1 ;
        RECT  0.000 0.000 0.620 234.760 ;
        LAYER metal2 ;
        RECT  0.000 0.000 0.620 234.760 ;
        LAYER metal3 ;
        RECT  0.000 0.000 0.620 234.760 ;
        LAYER metal4 ;
        RECT  0.000 0.000 0.620 234.760 ;
        LAYER metal5 ;
        RECT  0.000 0.000 0.620 234.760 ;
        LAYER metal6 ;
        RECT  0.000 0.000 0.620 234.760 ;
    END
END EMPTY1C

MACRO EMPTY1D
    CLASS PAD SPACER ;
    FOREIGN EMPTY1D 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.620 BY 140.120 ;
    SYMMETRY x y r90 ;
    SITE iocore_d ;
    OBS
        LAYER metal1 ;
        RECT  0.000 0.000 0.620 139.280 ;
        LAYER metal2 ;
        RECT  0.000 0.000 0.620 139.280 ;
        LAYER metal3 ;
        RECT  0.000 0.000 0.620 139.280 ;
        LAYER metal4 ;
        RECT  0.000 0.000 0.620 139.280 ;
        LAYER metal5 ;
        RECT  0.000 0.000 0.620 139.280 ;
        LAYER metal6 ;
        RECT  0.000 0.000 0.620 139.280 ;
    END
END EMPTY1D

MACRO EMPTY2C
    CLASS PAD SPACER ;
    FOREIGN EMPTY2C 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.240 BY 235.600 ;
    SYMMETRY x y r90 ;
    SITE iocore_c ;
    OBS
        LAYER metal1 ;
        RECT  0.000 0.000 1.240 234.760 ;
        LAYER metal2 ;
        RECT  0.000 0.000 1.240 234.760 ;
        LAYER metal3 ;
        RECT  0.000 0.000 1.240 234.760 ;
        LAYER metal4 ;
        RECT  0.000 0.000 1.240 234.760 ;
        LAYER metal5 ;
        RECT  0.000 0.000 1.240 234.760 ;
        LAYER metal6 ;
        RECT  0.000 0.000 1.240 234.760 ;
    END
END EMPTY2C

MACRO EMPTY2D
    CLASS PAD SPACER ;
    FOREIGN EMPTY2D 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.240 BY 140.120 ;
    SYMMETRY x y r90 ;
    SITE iocore_d ;
    OBS
        LAYER metal1 ;
        RECT  0.000 0.000 1.240 139.280 ;
        LAYER metal2 ;
        RECT  0.000 0.000 1.240 139.280 ;
        LAYER metal3 ;
        RECT  0.000 0.000 1.240 139.280 ;
        LAYER metal4 ;
        RECT  0.000 0.000 1.240 139.280 ;
        LAYER metal5 ;
        RECT  0.000 0.000 1.240 139.280 ;
        LAYER metal6 ;
        RECT  0.000 0.000 1.240 139.280 ;
    END
END EMPTY2D

MACRO EMPTY4C
    CLASS PAD SPACER ;
    FOREIGN EMPTY4C 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.480 BY 235.600 ;
    SYMMETRY x y r90 ;
    SITE iocore_c ;
    OBS
        LAYER metal1 ;
        RECT  0.000 0.000 2.480 234.760 ;
        LAYER metal2 ;
        RECT  0.000 0.000 2.480 234.760 ;
        LAYER metal3 ;
        RECT  0.000 0.000 2.480 234.760 ;
        LAYER metal4 ;
        RECT  0.000 0.000 2.480 234.760 ;
        LAYER metal5 ;
        RECT  0.000 0.000 2.480 234.760 ;
        LAYER metal6 ;
        RECT  0.000 0.000 2.480 234.760 ;
    END
END EMPTY4C

MACRO EMPTY4D
    CLASS PAD SPACER ;
    FOREIGN EMPTY4D 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.480 BY 140.120 ;
    SYMMETRY x y r90 ;
    SITE iocore_d ;
    OBS
        LAYER metal1 ;
        RECT  0.000 0.000 2.480 139.280 ;
        LAYER metal2 ;
        RECT  0.000 0.000 2.480 139.280 ;
        LAYER metal3 ;
        RECT  0.000 0.000 2.480 139.280 ;
        LAYER metal4 ;
        RECT  0.000 0.000 2.480 139.280 ;
        LAYER metal5 ;
        RECT  0.000 0.000 2.480 139.280 ;
        LAYER metal6 ;
        RECT  0.000 0.000 2.480 139.280 ;
    END
END EMPTY4D

MACRO EMPTY8C
    CLASS PAD SPACER ;
    FOREIGN EMPTY8C 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.960 BY 235.600 ;
    SYMMETRY x y r90 ;
    SITE iocore_c ;
    OBS
        LAYER metal1 ;
        RECT  0.000 0.000 4.960 234.760 ;
        LAYER metal2 ;
        RECT  0.000 0.000 4.960 234.760 ;
        LAYER metal3 ;
        RECT  0.000 0.000 4.960 234.760 ;
        LAYER metal4 ;
        RECT  0.000 0.000 4.960 234.760 ;
        LAYER metal5 ;
        RECT  0.000 0.000 4.960 234.760 ;
        LAYER metal6 ;
        RECT  0.000 0.000 4.960 234.760 ;
    END
END EMPTY8C

MACRO EMPTY8D
    CLASS PAD SPACER ;
    FOREIGN EMPTY8D 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.960 BY 140.120 ;
    SYMMETRY x y r90 ;
    SITE iocore_d ;
    OBS
        LAYER metal1 ;
        RECT  0.000 0.000 4.960 139.280 ;
        LAYER metal2 ;
        RECT  0.000 0.000 4.960 139.280 ;
        LAYER metal3 ;
        RECT  0.000 0.000 4.960 139.280 ;
        LAYER metal4 ;
        RECT  0.000 0.000 4.960 139.280 ;
        LAYER metal5 ;
        RECT  0.000 0.000 4.960 139.280 ;
        LAYER metal6 ;
        RECT  0.000 0.000 4.960 139.280 ;
    END
END EMPTY8D

MACRO EMPTYGRC
    CLASS PAD SPACER ;
    FOREIGN EMPTYGRC 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.720 BY 235.600 ;
    SYMMETRY x y r90 ;
    SITE iocore_c ;
    OBS
        LAYER metal1 ;
        RECT  0.000 0.000 3.720 234.760 ;
        LAYER metal2 ;
        RECT  0.000 0.000 3.720 234.760 ;
        LAYER metal3 ;
        RECT  0.000 0.000 3.720 234.760 ;
        LAYER metal4 ;
        RECT  0.000 0.000 3.720 234.760 ;
        LAYER metal5 ;
        RECT  0.000 0.000 3.720 234.760 ;
        LAYER metal6 ;
        RECT  0.000 0.000 3.720 234.760 ;
    END
END EMPTYGRC

MACRO EMPTYGRD
    CLASS PAD SPACER ;
    FOREIGN EMPTYGRD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.720 BY 140.120 ;
    SYMMETRY x y r90 ;
    SITE iocore_d ;
    OBS
        LAYER metal1 ;
        RECT  0.000 0.000 3.720 139.280 ;
        LAYER metal2 ;
        RECT  0.000 0.000 3.720 139.280 ;
        LAYER metal3 ;
        RECT  0.000 0.000 3.720 139.280 ;
        LAYER metal4 ;
        RECT  0.000 0.000 3.720 139.280 ;
        LAYER metal5 ;
        RECT  0.000 0.000 3.720 139.280 ;
        LAYER metal6 ;
        RECT  0.000 0.000 3.720 139.280 ;
    END
END EMPTYGRD

MACRO GNDIOC
    CLASS PAD ;
    FOREIGN GNDIOC 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 34.100 BY 235.600 ;
    SYMMETRY x y r90 ;
    SITE iocore_c ;
    PIN GNDO
        DIRECTION INOUT ;
        USE ANALOG ;
        PORT
        LAYER metal6 ;
        RECT  1.910 0.000 32.190 4.300 ;
        LAYER metal5 ;
        RECT  1.910 0.000 32.190 4.300 ;
        LAYER metal4 ;
        RECT  1.910 0.000 32.190 4.300 ;
        LAYER metal3 ;
        RECT  1.910 0.000 32.190 4.300 ;
        LAYER metal2 ;
        RECT  1.910 0.000 32.190 4.300 ;
        LAYER metal1 ;
        RECT  1.910 0.000 32.190 4.300 ;
        END
    END GNDO
    OBS
        LAYER metal1 ;
        POLYGON  34.100 235.600 0.000 235.600 0.000 0.000 1.630 0.000 1.630 4.580
                 32.470 4.580 32.470 0.000 34.100 0.000 ;
        LAYER via ;
        RECT  1.910 0.000 32.190 4.300 ;
        LAYER metal2 ;
        POLYGON  34.100 235.600 0.000 235.600 0.000 0.000 1.590 0.000 1.590 4.620
                 32.510 4.620 32.510 0.000 34.100 0.000 ;
        LAYER via2 ;
        RECT  1.910 0.000 32.190 4.300 ;
        LAYER metal3 ;
        POLYGON  34.100 235.600 0.000 235.600 0.000 0.000 1.590 0.000 1.590 4.620
                 32.510 4.620 32.510 0.000 34.100 0.000 ;
        LAYER via3 ;
        RECT  1.910 0.000 32.190 4.300 ;
        LAYER metal4 ;
        POLYGON  34.100 235.600 0.000 235.600 0.000 0.000 1.590 0.000 1.590 4.620
                 32.510 4.620 32.510 0.000 34.100 0.000 ;
        LAYER via4 ;
        RECT  1.910 0.000 32.190 4.300 ;
        LAYER metal5 ;
        POLYGON  34.100 235.600 0.000 235.600 0.000 0.000 1.590 0.000 1.590 4.620
                 32.510 4.620 32.510 0.000 34.100 0.000 ;
        LAYER via5 ;
        RECT  1.910 0.000 32.190 4.300 ;
        LAYER metal6 ;
        POLYGON  34.100 235.600 0.000 235.600 0.000 0.000 1.310 0.000 1.310 4.900
                 32.790 4.900 32.790 0.000 34.100 0.000 ;
    END
END GNDIOC

MACRO GNDIOD
    CLASS PAD ;
    FOREIGN GNDIOD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 62.620 BY 140.120 ;
    SYMMETRY x y r90 ;
    SITE iocore_d ;
    PIN GNDO
        DIRECTION INOUT ;
        USE ANALOG ;
        PORT
        LAYER metal6 ;
        RECT  2.850 0.000 59.770 3.000 ;
        LAYER metal5 ;
        RECT  2.850 0.000 59.770 3.000 ;
        LAYER metal4 ;
        RECT  2.850 0.000 59.770 3.000 ;
        LAYER metal3 ;
        RECT  2.850 0.000 59.770 3.000 ;
        LAYER metal2 ;
        RECT  2.850 0.000 59.770 3.000 ;
        LAYER metal1 ;
        RECT  2.850 0.000 59.770 3.000 ;
        END
    END GNDO
    OBS
        LAYER metal1 ;
        POLYGON  62.620 140.120 0.000 140.120 0.000 0.000 2.570 0.000 2.570 3.280
                 60.050 3.280 60.050 0.000 62.620 0.000 ;
        LAYER via ;
        RECT  2.850 0.000 59.770 3.000 ;
        LAYER metal2 ;
        POLYGON  62.620 140.120 0.000 140.120 0.000 0.000 2.530 0.000 2.530 3.320
                 60.090 3.320 60.090 0.000 62.620 0.000 ;
        LAYER via2 ;
        RECT  2.850 0.000 59.770 3.000 ;
        LAYER metal3 ;
        POLYGON  62.620 140.120 0.000 140.120 0.000 0.000 2.530 0.000 2.530 3.320
                 60.090 3.320 60.090 0.000 62.620 0.000 ;
        LAYER via3 ;
        RECT  2.850 0.000 59.770 3.000 ;
        LAYER metal4 ;
        POLYGON  62.620 140.120 0.000 140.120 0.000 0.000 2.530 0.000 2.530 3.320
                 60.090 3.320 60.090 0.000 62.620 0.000 ;
        LAYER via4 ;
        RECT  2.850 0.000 59.770 3.000 ;
        LAYER metal5 ;
        POLYGON  62.620 140.120 0.000 140.120 0.000 0.000 2.530 0.000 2.530 3.320
                 60.090 3.320 60.090 0.000 62.620 0.000 ;
        LAYER via5 ;
        RECT  2.850 0.000 59.770 3.000 ;
        LAYER metal6 ;
        POLYGON  62.620 140.120 0.000 140.120 0.000 0.000 2.250 0.000 2.250 3.600
                 60.370 3.600 60.370 0.000 62.620 0.000 ;
    END
END GNDIOD

MACRO GNDKC
    CLASS PAD ;
    FOREIGN GNDKC 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 34.100 BY 235.600 ;
    SYMMETRY x y r90 ;
    SITE iocore_c ;
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        PORT
        CLASS CORE ;
        LAYER metal6 ;
        RECT  18.050 231.090 32.090 235.360 ;
        LAYER metal5 ;
        RECT  18.050 231.090 32.090 235.360 ;
        LAYER metal4 ;
        RECT  18.050 231.090 32.090 235.360 ;
        LAYER metal3 ;
        RECT  18.050 231.090 32.090 235.360 ;
        LAYER metal2 ;
        RECT  18.050 231.090 32.090 235.360 ;
        LAYER metal1 ;
        RECT  18.050 231.090 32.090 235.360 ;
        END
        PORT
        CLASS CORE ;
        LAYER metal6 ;
        RECT  2.010 231.090 16.050 235.360 ;
        LAYER metal5 ;
        RECT  2.010 231.090 16.050 235.360 ;
        LAYER metal4 ;
        RECT  2.010 231.090 16.050 235.360 ;
        LAYER metal3 ;
        RECT  2.010 231.090 16.050 235.360 ;
        LAYER metal2 ;
        RECT  2.010 231.090 16.050 235.360 ;
        LAYER metal1 ;
        RECT  2.010 231.090 16.050 235.360 ;
        END
        PORT
        CLASS CORE ;
        LAYER metal6 ;
        RECT  1.910 0.000 32.190 4.300 ;
        LAYER metal5 ;
        RECT  1.910 0.000 32.190 4.300 ;
        LAYER metal4 ;
        RECT  1.910 0.000 32.190 4.300 ;
        LAYER metal3 ;
        RECT  1.910 0.000 32.190 4.300 ;
        LAYER metal2 ;
        RECT  1.910 0.000 32.190 4.300 ;
        LAYER metal1 ;
        RECT  1.910 0.000 32.190 4.300 ;
        END
    END GND
    OBS
        LAYER metal1 ;
        POLYGON  34.100 235.360 32.370 235.360 32.370 230.810 17.770 230.810
                 17.770 235.360 16.330 235.360 16.330 230.810 1.730 230.810 1.730 235.360
                 0.000 235.360 0.000 0.000 1.630 0.000 1.630 4.580 32.470 4.580
                 32.470 0.000 34.100 0.000 ;
        LAYER via ;
        RECT  18.050 231.090 32.090 235.360 ;
        RECT  2.010 231.090 16.050 235.360 ;
        RECT  1.910 0.000 32.190 4.300 ;
        LAYER metal2 ;
        POLYGON  34.100 235.360 32.410 235.360 32.410 230.770 17.730 230.770
                 17.730 235.360 16.370 235.360 16.370 230.770 1.690 230.770 1.690 235.360
                 0.000 235.360 0.000 0.000 1.590 0.000 1.590 4.620 32.510 4.620
                 32.510 0.000 34.100 0.000 ;
        LAYER via2 ;
        RECT  18.050 231.090 32.090 235.360 ;
        RECT  2.010 231.090 16.050 235.360 ;
        RECT  1.910 0.000 32.190 4.300 ;
        LAYER metal3 ;
        POLYGON  34.100 235.360 32.410 235.360 32.410 230.770 17.730 230.770
                 17.730 235.360 16.370 235.360 16.370 230.770 1.690 230.770 1.690 235.360
                 0.000 235.360 0.000 0.000 1.590 0.000 1.590 4.620 32.510 4.620
                 32.510 0.000 34.100 0.000 ;
        LAYER via3 ;
        RECT  18.050 231.090 32.090 235.360 ;
        RECT  2.010 231.090 16.050 235.360 ;
        RECT  1.910 0.000 32.190 4.300 ;
        LAYER metal4 ;
        POLYGON  34.100 235.360 32.410 235.360 32.410 230.770 17.730 230.770
                 17.730 235.360 16.370 235.360 16.370 230.770 1.690 230.770 1.690 235.360
                 0.000 235.360 0.000 0.000 1.590 0.000 1.590 4.620 32.510 4.620
                 32.510 0.000 34.100 0.000 ;
        LAYER via4 ;
        RECT  18.050 231.090 32.090 235.360 ;
        RECT  2.010 231.090 16.050 235.360 ;
        RECT  1.910 0.000 32.190 4.300 ;
        LAYER metal5 ;
        POLYGON  34.100 235.360 32.410 235.360 32.410 230.770 17.730 230.770
                 17.730 235.360 16.370 235.360 16.370 230.770 1.690 230.770 1.690 235.360
                 0.000 235.360 0.000 0.000 1.590 0.000 1.590 4.620 32.510 4.620
                 32.510 0.000 34.100 0.000 ;
        LAYER via5 ;
        RECT  18.050 231.090 32.090 235.360 ;
        RECT  2.010 231.090 16.050 235.360 ;
        RECT  1.910 0.000 32.190 4.300 ;
        LAYER metal6 ;
        POLYGON  34.100 235.360 32.690 235.360 32.690 230.490 17.450 230.490
                 17.450 235.360 16.650 235.360 16.650 230.490 1.410 230.490 1.410 235.360
                 0.000 235.360 0.000 0.000 1.310 0.000 1.310 4.900 32.790 4.900
                 32.790 0.000 34.100 0.000 ;
    END
END GNDKC

MACRO GNDKD
    CLASS PAD ;
    FOREIGN GNDKD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 62.620 BY 140.120 ;
    SYMMETRY x y r90 ;
    SITE iocore_d ;
    PIN GND
        DIRECTION INOUT ;
        USE ground ;
        PORT
        CLASS CORE ;
        LAYER metal6 ;
        RECT  2.850 0.000 59.770 3.000 ;
        LAYER metal5 ;
        RECT  2.850 0.000 59.770 3.000 ;
        LAYER metal4 ;
        RECT  2.850 0.000 59.770 3.000 ;
        LAYER metal3 ;
        RECT  2.850 0.000 59.770 3.000 ;
        LAYER metal2 ;
        RECT  2.850 0.000 59.770 3.000 ;
        LAYER metal1 ;
        RECT  2.850 0.000 59.770 3.000 ;
        END
        PORT
        CLASS CORE ;
        LAYER metal6 ;
        RECT  42.310 135.360 60.210 139.880 ;
        LAYER metal5 ;
        RECT  42.310 135.360 60.210 139.880 ;
        LAYER metal4 ;
        RECT  42.310 135.360 60.210 139.880 ;
        LAYER metal3 ;
        RECT  42.310 135.360 60.210 139.880 ;
        LAYER metal2 ;
        RECT  42.310 135.360 60.210 139.880 ;
        LAYER metal1 ;
        RECT  42.310 135.360 60.210 139.880 ;
        END
        PORT
        CLASS CORE ;
        LAYER metal6 ;
        RECT  22.310 135.360 40.310 139.880 ;
        LAYER metal5 ;
        RECT  22.310 135.360 40.310 139.880 ;
        LAYER metal4 ;
        RECT  22.310 135.360 40.310 139.880 ;
        LAYER metal3 ;
        RECT  22.310 135.360 40.310 139.880 ;
        LAYER metal2 ;
        RECT  22.310 135.360 40.310 139.880 ;
        LAYER metal1 ;
        RECT  22.310 135.360 40.310 139.880 ;
        END
        PORT
        CLASS CORE ;
        LAYER metal6 ;
        RECT  2.410 135.360 20.310 139.880 ;
        LAYER metal5 ;
        RECT  2.410 135.360 20.310 139.880 ;
        LAYER metal4 ;
        RECT  2.410 135.360 20.310 139.880 ;
        LAYER metal3 ;
        RECT  2.410 135.360 20.310 139.880 ;
        LAYER metal2 ;
        RECT  2.410 135.360 20.310 139.880 ;
        LAYER metal1 ;
        RECT  2.410 135.360 20.310 139.880 ;
        END
    END GND
    OBS
        LAYER metal1 ;
        POLYGON  62.620 139.880 60.490 139.880 60.490 135.080 42.030 135.080
                 42.030 139.880 40.590 139.880 40.590 135.080 22.030 135.080
                 22.030 139.880 20.590 139.880 20.590 135.080 2.130 135.080 2.130 139.880
                 0.000 139.880 0.000 0.000 2.570 0.000 2.570 3.280 60.050 3.280
                 60.050 0.000 62.620 0.000 ;
        LAYER via ;
        RECT  2.850 0.000 59.770 3.000 ;
        RECT  42.310 135.360 60.210 139.880 ;
        RECT  22.310 135.360 40.310 139.880 ;
        RECT  2.410 135.360 20.310 139.880 ;
        LAYER metal2 ;
        POLYGON  62.620 139.880 60.530 139.880 60.530 135.040 41.990 135.040
                 41.990 139.880 40.630 139.880 40.630 135.040 21.990 135.040
                 21.990 139.880 20.630 139.880 20.630 135.040 2.090 135.040 2.090 139.880
                 0.000 139.880 0.000 0.000 2.530 0.000 2.530 3.320 60.090 3.320
                 60.090 0.000 62.620 0.000 ;
        LAYER via2 ;
        RECT  2.850 0.000 59.770 3.000 ;
        RECT  42.310 135.360 60.210 139.880 ;
        RECT  22.310 135.360 40.310 139.880 ;
        RECT  2.410 135.360 20.310 139.880 ;
        LAYER metal3 ;
        POLYGON  62.620 139.880 60.530 139.880 60.530 135.040 41.990 135.040
                 41.990 139.880 40.630 139.880 40.630 135.040 21.990 135.040
                 21.990 139.880 20.630 139.880 20.630 135.040 2.090 135.040 2.090 139.880
                 0.000 139.880 0.000 0.000 2.530 0.000 2.530 3.320 60.090 3.320
                 60.090 0.000 62.620 0.000 ;
        LAYER via3 ;
        RECT  2.850 0.000 59.770 3.000 ;
        RECT  42.310 135.360 60.210 139.880 ;
        RECT  22.310 135.360 40.310 139.880 ;
        RECT  2.410 135.360 20.310 139.880 ;
        LAYER metal4 ;
        POLYGON  62.620 139.880 60.530 139.880 60.530 135.040 41.990 135.040
                 41.990 139.880 40.630 139.880 40.630 135.040 21.990 135.040
                 21.990 139.880 20.630 139.880 20.630 135.040 2.090 135.040 2.090 139.880
                 0.000 139.880 0.000 0.000 2.530 0.000 2.530 3.320 60.090 3.320
                 60.090 0.000 62.620 0.000 ;
        LAYER via4 ;
        RECT  2.850 0.000 59.770 3.000 ;
        RECT  42.310 135.360 60.210 139.880 ;
        RECT  22.310 135.360 40.310 139.880 ;
        RECT  2.410 135.360 20.310 139.880 ;
        LAYER metal5 ;
        POLYGON  62.620 139.880 60.530 139.880 60.530 135.040 41.990 135.040
                 41.990 139.880 40.630 139.880 40.630 135.040 21.990 135.040
                 21.990 139.880 20.630 139.880 20.630 135.040 2.090 135.040 2.090 139.880
                 0.000 139.880 0.000 0.000 2.530 0.000 2.530 3.320 60.090 3.320
                 60.090 0.000 62.620 0.000 ;
        LAYER via5 ;
        RECT  2.850 0.000 59.770 3.000 ;
        RECT  42.310 135.360 60.210 139.880 ;
        RECT  22.310 135.360 40.310 139.880 ;
        RECT  2.410 135.360 20.310 139.880 ;
        LAYER metal6 ;
        POLYGON  62.620 139.880 60.810 139.880 60.810 134.760 41.710 134.760
                 41.710 139.880 40.910 139.880 40.910 134.760 21.710 134.760
                 21.710 139.880 20.910 139.880 20.910 134.760 1.810 134.760 1.810 139.880
                 0.000 139.880 0.000 0.000 2.250 0.000 2.250 3.600 60.370 3.600
                 60.370 0.000 62.620 0.000 ;
    END
END GNDKD

MACRO VCC3IOC
    CLASS PAD ;
    FOREIGN VCC3IOC 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 34.100 BY 235.600 ;
    SYMMETRY x y r90 ;
    SITE iocore_c ;
    PIN VCC3O
        DIRECTION INOUT ;
        USE ANALOG ;
        PORT
        LAYER metal6 ;
        RECT  1.910 0.000 32.190 4.300 ;
        LAYER metal5 ;
        RECT  1.910 0.000 32.190 4.300 ;
        LAYER metal4 ;
        RECT  1.910 0.000 32.190 4.300 ;
        LAYER metal3 ;
        RECT  1.910 0.000 32.190 4.300 ;
        LAYER metal2 ;
        RECT  1.910 0.000 32.190 4.300 ;
        LAYER metal1 ;
        RECT  1.910 0.000 32.190 4.300 ;
        END
    END VCC3O
    OBS
        LAYER metal1 ;
        POLYGON  34.100 235.600 0.000 235.600 0.000 0.000 1.630 0.000 1.630 4.580
                 32.470 4.580 32.470 0.000 34.100 0.000 ;
        LAYER via ;
        RECT  1.910 0.000 32.190 4.300 ;
        LAYER metal2 ;
        POLYGON  34.100 235.600 0.000 235.600 0.000 0.000 1.590 0.000 1.590 4.620
                 32.510 4.620 32.510 0.000 34.100 0.000 ;
        LAYER via2 ;
        RECT  1.910 0.000 32.190 4.300 ;
        LAYER metal3 ;
        POLYGON  34.100 235.600 0.000 235.600 0.000 0.000 1.590 0.000 1.590 4.620
                 32.510 4.620 32.510 0.000 34.100 0.000 ;
        LAYER via3 ;
        RECT  1.910 0.000 32.190 4.300 ;
        LAYER metal4 ;
        POLYGON  34.100 235.600 0.000 235.600 0.000 0.000 1.590 0.000 1.590 4.620
                 32.510 4.620 32.510 0.000 34.100 0.000 ;
        LAYER via4 ;
        RECT  1.910 0.000 32.190 4.300 ;
        LAYER metal5 ;
        POLYGON  34.100 235.600 0.000 235.600 0.000 0.000 1.590 0.000 1.590 4.620
                 32.510 4.620 32.510 0.000 34.100 0.000 ;
        LAYER via5 ;
        RECT  1.910 0.000 32.190 4.300 ;
        LAYER metal6 ;
        POLYGON  34.100 235.600 0.000 235.600 0.000 0.000 1.310 0.000 1.310 4.900
                 32.790 4.900 32.790 0.000 34.100 0.000 ;
    END
END VCC3IOC

MACRO VCC3IOD
    CLASS PAD ;
    FOREIGN VCC3IOD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 62.620 BY 140.120 ;
    SYMMETRY x y r90 ;
    SITE iocore_d ;
    PIN VCC3O
        DIRECTION INOUT ;
        USE ANALOG ;
        PORT
        LAYER metal6 ;
        RECT  2.850 0.000 59.770 3.000 ;
        LAYER metal5 ;
        RECT  2.850 0.000 59.770 3.000 ;
        LAYER metal4 ;
        RECT  2.850 0.000 59.770 3.000 ;
        LAYER metal3 ;
        RECT  2.850 0.000 59.770 3.000 ;
        LAYER metal2 ;
        RECT  2.850 0.000 59.770 3.000 ;
        LAYER metal1 ;
        RECT  2.850 0.000 59.770 3.000 ;
        END
    END VCC3O
    OBS
        LAYER metal1 ;
        POLYGON  62.620 140.120 0.000 140.120 0.000 0.000 2.570 0.000 2.570 3.280
                 60.050 3.280 60.050 0.000 62.620 0.000 ;
        LAYER via ;
        RECT  2.850 0.000 59.770 3.000 ;
        LAYER metal2 ;
        POLYGON  62.620 140.120 0.000 140.120 0.000 0.000 2.530 0.000 2.530 3.320
                 60.090 3.320 60.090 0.000 62.620 0.000 ;
        LAYER via2 ;
        RECT  2.850 0.000 59.770 3.000 ;
        LAYER metal3 ;
        POLYGON  62.620 140.120 0.000 140.120 0.000 0.000 2.530 0.000 2.530 3.320
                 60.090 3.320 60.090 0.000 62.620 0.000 ;
        LAYER via3 ;
        RECT  2.850 0.000 59.770 3.000 ;
        LAYER metal4 ;
        POLYGON  62.620 140.120 0.000 140.120 0.000 0.000 2.530 0.000 2.530 3.320
                 60.090 3.320 60.090 0.000 62.620 0.000 ;
        LAYER via4 ;
        RECT  2.850 0.000 59.770 3.000 ;
        LAYER metal5 ;
        POLYGON  62.620 140.120 0.000 140.120 0.000 0.000 2.530 0.000 2.530 3.320
                 60.090 3.320 60.090 0.000 62.620 0.000 ;
        LAYER via5 ;
        RECT  2.850 0.000 59.770 3.000 ;
        LAYER metal6 ;
        POLYGON  62.620 140.120 0.000 140.120 0.000 0.000 2.250 0.000 2.250 3.600
                 60.370 3.600 60.370 0.000 62.620 0.000 ;
    END
END VCC3IOD

MACRO VCCKC
    CLASS PAD ;
    FOREIGN VCCKC 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 34.100 BY 235.600 ;
    SYMMETRY x y r90 ;
    SITE iocore_c ;
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        PORT
        CLASS CORE ;
        LAYER metal6 ;
        RECT  1.910 0.000 32.190 4.300 ;
        LAYER metal5 ;
        RECT  1.910 0.000 32.190 4.300 ;
        LAYER metal4 ;
        RECT  1.910 0.000 32.190 4.300 ;
        LAYER metal3 ;
        RECT  1.910 0.000 32.190 4.300 ;
        LAYER metal2 ;
        RECT  1.910 0.000 32.190 4.300 ;
        LAYER metal1 ;
        RECT  1.910 0.000 32.190 4.300 ;
        END
        PORT
        CLASS CORE ;
        LAYER metal6 ;
        RECT  18.050 231.090 32.190 235.360 ;
        LAYER metal5 ;
        RECT  18.050 231.090 32.190 235.360 ;
        LAYER metal4 ;
        RECT  18.050 231.090 32.190 235.360 ;
        LAYER metal3 ;
        RECT  18.050 231.090 32.190 235.360 ;
        LAYER metal2 ;
        RECT  18.050 231.090 32.190 235.360 ;
        LAYER metal1 ;
        RECT  18.050 231.090 32.190 235.360 ;
        END
        PORT
        CLASS CORE ;
        LAYER metal6 ;
        RECT  1.910 231.090 16.050 235.360 ;
        LAYER metal5 ;
        RECT  1.910 231.090 16.050 235.360 ;
        LAYER metal4 ;
        RECT  1.910 231.090 16.050 235.360 ;
        LAYER metal3 ;
        RECT  1.910 231.090 16.050 235.360 ;
        LAYER metal2 ;
        RECT  1.910 231.090 16.050 235.360 ;
        LAYER metal1 ;
        RECT  1.910 231.090 16.050 235.360 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        POLYGON  34.100 235.360 32.470 235.360 32.470 230.810 17.770 230.810
                 17.770 235.360 16.330 235.360 16.330 230.810 1.630 230.810 1.630 235.360
                 0.000 235.360 0.000 0.000 1.630 0.000 1.630 4.580 32.470 4.580
                 32.470 0.000 34.100 0.000 ;
        LAYER via ;
        RECT  1.910 0.000 32.190 4.300 ;
        RECT  18.050 231.090 32.190 235.360 ;
        RECT  1.910 231.090 16.050 235.360 ;
        LAYER metal2 ;
        POLYGON  34.100 235.360 32.510 235.360 32.510 230.770 17.730 230.770
                 17.730 235.360 16.370 235.360 16.370 230.770 1.590 230.770 1.590 235.360
                 0.000 235.360 0.000 0.000 1.590 0.000 1.590 4.620 32.510 4.620
                 32.510 0.000 34.100 0.000 ;
        LAYER via2 ;
        RECT  1.910 0.000 32.190 4.300 ;
        RECT  18.050 231.090 32.190 235.360 ;
        RECT  1.910 231.090 16.050 235.360 ;
        LAYER metal3 ;
        POLYGON  34.100 235.360 32.510 235.360 32.510 230.770 17.730 230.770
                 17.730 235.360 16.370 235.360 16.370 230.770 1.590 230.770 1.590 235.360
                 0.000 235.360 0.000 0.000 1.590 0.000 1.590 4.620 32.510 4.620
                 32.510 0.000 34.100 0.000 ;
        LAYER via3 ;
        RECT  1.910 0.000 32.190 4.300 ;
        RECT  18.050 231.090 32.190 235.360 ;
        RECT  1.910 231.090 16.050 235.360 ;
        LAYER metal4 ;
        POLYGON  34.100 235.360 32.510 235.360 32.510 230.770 17.730 230.770
                 17.730 235.360 16.370 235.360 16.370 230.770 1.590 230.770 1.590 235.360
                 0.000 235.360 0.000 0.000 1.590 0.000 1.590 4.620 32.510 4.620
                 32.510 0.000 34.100 0.000 ;
        LAYER via4 ;
        RECT  1.910 0.000 32.190 4.300 ;
        RECT  18.050 231.090 32.190 235.360 ;
        RECT  1.910 231.090 16.050 235.360 ;
        LAYER metal5 ;
        POLYGON  34.100 235.360 32.510 235.360 32.510 230.770 17.730 230.770
                 17.730 235.360 16.370 235.360 16.370 230.770 1.590 230.770 1.590 235.360
                 0.000 235.360 0.000 0.000 1.590 0.000 1.590 4.620 32.510 4.620
                 32.510 0.000 34.100 0.000 ;
        LAYER via5 ;
        RECT  1.910 0.000 32.190 4.300 ;
        RECT  18.050 231.090 32.190 235.360 ;
        RECT  1.910 231.090 16.050 235.360 ;
        LAYER metal6 ;
        POLYGON  34.100 235.360 32.790 235.360 32.790 230.490 17.450 230.490
                 17.450 235.360 16.650 235.360 16.650 230.490 1.310 230.490 1.310 235.360
                 0.000 235.360 0.000 0.000 1.310 0.000 1.310 4.900 32.790 4.900
                 32.790 0.000 34.100 0.000 ;
    END
END VCCKC

MACRO VCCKD
    CLASS PAD ;
    FOREIGN VCCKD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 62.620 BY 140.120 ;
    SYMMETRY x y r90 ;
    SITE iocore_d ;
    PIN VCC
        DIRECTION INOUT ;
        USE power ;
        PORT
        CLASS CORE ;
        LAYER metal6 ;
        RECT  2.850 0.000 59.770 3.000 ;
        LAYER metal5 ;
        RECT  2.850 0.000 59.770 3.000 ;
        LAYER metal4 ;
        RECT  2.850 0.000 59.770 3.000 ;
        LAYER metal3 ;
        RECT  2.850 0.000 59.770 3.000 ;
        LAYER metal2 ;
        RECT  2.850 0.000 59.770 3.000 ;
        LAYER metal1 ;
        RECT  2.850 0.000 59.770 3.000 ;
        END
        PORT
        CLASS CORE ;
        LAYER metal6 ;
        RECT  2.850 135.360 20.490 139.880 ;
        LAYER metal5 ;
        RECT  2.850 135.360 20.490 139.880 ;
        LAYER metal4 ;
        RECT  2.850 135.360 20.490 139.880 ;
        LAYER metal3 ;
        RECT  2.850 135.360 20.490 139.880 ;
        LAYER metal2 ;
        RECT  2.850 135.360 20.490 139.880 ;
        LAYER metal1 ;
        RECT  2.850 135.360 20.490 139.880 ;
        END
        PORT
        CLASS CORE ;
        LAYER metal6 ;
        RECT  22.490 135.360 40.130 139.880 ;
        LAYER metal5 ;
        RECT  22.490 135.360 40.130 139.880 ;
        LAYER metal4 ;
        RECT  22.490 135.360 40.130 139.880 ;
        LAYER metal3 ;
        RECT  22.490 135.360 40.130 139.880 ;
        LAYER metal2 ;
        RECT  22.490 135.360 40.130 139.880 ;
        LAYER metal1 ;
        RECT  22.490 135.360 40.130 139.880 ;
        END
        PORT
        CLASS CORE ;
        LAYER metal6 ;
        RECT  42.130 135.360 59.770 139.880 ;
        LAYER metal5 ;
        RECT  42.130 135.360 59.770 139.880 ;
        LAYER metal4 ;
        RECT  42.130 135.360 59.770 139.880 ;
        LAYER metal3 ;
        RECT  42.130 135.360 59.770 139.880 ;
        LAYER metal2 ;
        RECT  42.130 135.360 59.770 139.880 ;
        LAYER metal1 ;
        RECT  42.130 135.360 59.770 139.880 ;
        END
    END VCC
    OBS
        LAYER metal1 ;
        POLYGON  62.620 139.880 60.050 139.880 60.050 135.080 41.850 135.080
                 41.850 139.880 40.410 139.880 40.410 135.080 22.210 135.080
                 22.210 139.880 20.770 139.880 20.770 135.080 2.570 135.080 2.570 139.880
                 0.000 139.880 0.000 0.000 2.570 0.000 2.570 3.280 60.050 3.280
                 60.050 0.000 62.620 0.000 ;
        LAYER via ;
        RECT  2.850 0.000 59.770 3.000 ;
        RECT  2.850 135.360 20.490 139.880 ;
        RECT  22.490 135.360 40.130 139.880 ;
        RECT  42.130 135.360 59.770 139.880 ;
        LAYER metal2 ;
        POLYGON  62.620 139.880 60.090 139.880 60.090 135.040 41.810 135.040
                 41.810 139.880 40.450 139.880 40.450 135.040 22.170 135.040
                 22.170 139.880 20.810 139.880 20.810 135.040 2.530 135.040 2.530 139.880
                 0.000 139.880 0.000 0.000 2.530 0.000 2.530 3.320 60.090 3.320
                 60.090 0.000 62.620 0.000 ;
        LAYER via2 ;
        RECT  2.850 0.000 59.770 3.000 ;
        RECT  2.850 135.360 20.490 139.880 ;
        RECT  22.490 135.360 40.130 139.880 ;
        RECT  42.130 135.360 59.770 139.880 ;
        LAYER metal3 ;
        POLYGON  62.620 139.880 60.090 139.880 60.090 135.040 41.810 135.040
                 41.810 139.880 40.450 139.880 40.450 135.040 22.170 135.040
                 22.170 139.880 20.810 139.880 20.810 135.040 2.530 135.040 2.530 139.880
                 0.000 139.880 0.000 0.000 2.530 0.000 2.530 3.320 60.090 3.320
                 60.090 0.000 62.620 0.000 ;
        LAYER via3 ;
        RECT  2.850 0.000 59.770 3.000 ;
        RECT  2.850 135.360 20.490 139.880 ;
        RECT  22.490 135.360 40.130 139.880 ;
        RECT  42.130 135.360 59.770 139.880 ;
        LAYER metal4 ;
        POLYGON  62.620 139.880 60.090 139.880 60.090 135.040 41.810 135.040
                 41.810 139.880 40.450 139.880 40.450 135.040 22.170 135.040
                 22.170 139.880 20.810 139.880 20.810 135.040 2.530 135.040 2.530 139.880
                 0.000 139.880 0.000 0.000 2.530 0.000 2.530 3.320 60.090 3.320
                 60.090 0.000 62.620 0.000 ;
        LAYER via4 ;
        RECT  2.850 0.000 59.770 3.000 ;
        RECT  2.850 135.360 20.490 139.880 ;
        RECT  22.490 135.360 40.130 139.880 ;
        RECT  42.130 135.360 59.770 139.880 ;
        LAYER metal5 ;
        POLYGON  62.620 139.880 60.090 139.880 60.090 135.040 41.810 135.040
                 41.810 139.880 40.450 139.880 40.450 135.040 22.170 135.040
                 22.170 139.880 20.810 139.880 20.810 135.040 2.530 135.040 2.530 139.880
                 0.000 139.880 0.000 0.000 2.530 0.000 2.530 3.320 60.090 3.320
                 60.090 0.000 62.620 0.000 ;
        LAYER via5 ;
        RECT  2.850 0.000 59.770 3.000 ;
        RECT  2.850 135.360 20.490 139.880 ;
        RECT  22.490 135.360 40.130 139.880 ;
        RECT  42.130 135.360 59.770 139.880 ;
        LAYER metal6 ;
        POLYGON  62.620 139.880 60.370 139.880 60.370 134.760 41.530 134.760
                 41.530 139.880 40.730 139.880 40.730 134.760 21.890 134.760
                 21.890 139.880 21.090 139.880 21.090 134.760 2.250 134.760 2.250 139.880
                 0.000 139.880 0.000 0.000 2.250 0.000 2.250 3.600 60.370 3.600
                 60.370 0.000 62.620 0.000 ;
    END
END VCCKD

MACRO XMC
    CLASS PAD ;
    FOREIGN XMC 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 34.100 BY 235.600 ;
    SYMMETRY x y r90 ;
    SITE iocore_c ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal3 ;
        RECT  15.490 234.080 17.370 234.980 ;
        LAYER metal2 ;
        RECT  15.490 234.080 17.370 234.980 ;
        LAYER metal1 ;
        RECT  15.490 234.080 17.370 234.980 ;
        END
    END O
    PIN PD
        DIRECTION INPUT ;
        PORT
        LAYER metal3 ;
        RECT  9.290 234.080 11.170 234.980 ;
        LAYER metal2 ;
        RECT  9.290 234.080 11.170 234.980 ;
        LAYER metal1 ;
        RECT  9.290 234.080 11.170 234.980 ;
        END
    END PD
    PIN PU
        DIRECTION INPUT ;
        PORT
        LAYER metal3 ;
        RECT  5.570 234.080 7.450 234.980 ;
        LAYER metal2 ;
        RECT  5.570 234.080 7.450 234.980 ;
        LAYER metal1 ;
        RECT  5.570 234.080 7.450 234.980 ;
        END
    END PU
    PIN SMT
        DIRECTION INPUT ;
        PORT
        LAYER metal3 ;
        RECT  1.850 234.080 3.730 234.980 ;
        LAYER metal2 ;
        RECT  1.850 234.080 3.730 234.980 ;
        LAYER metal1 ;
        RECT  1.850 234.080 3.730 234.980 ;
        END
    END SMT
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal6 ;
        RECT  1.910 0.000 32.190 4.300 ;
        LAYER metal5 ;
        RECT  1.910 0.000 32.190 4.300 ;
        LAYER metal4 ;
        RECT  1.910 0.000 32.190 4.300 ;
        LAYER metal3 ;
        RECT  1.910 0.000 32.190 4.300 ;
        LAYER metal2 ;
        RECT  1.910 0.000 32.190 4.300 ;
        LAYER metal1 ;
        RECT  1.910 0.000 32.190 4.300 ;
        END
    END I
    OBS
        LAYER metal1 ;
        POLYGON  34.100 234.980 17.610 234.980 17.610 233.840 15.250 233.840
                 15.250 234.980 11.410 234.980 11.410 233.840 9.050 233.840 9.050 234.980
                 7.690 234.980 7.690 233.840 5.330 233.840 5.330 234.980 3.970 234.980
                 3.970 233.840 1.610 233.840 1.610 234.980 0.000 234.980 0.000 0.000
                 1.630 0.000 1.630 4.580 32.470 4.580 32.470 0.000 34.100 0.000 ;
        LAYER via ;
        RECT  15.490 234.080 17.370 234.980 ;
        RECT  9.290 234.080 11.170 234.980 ;
        RECT  5.570 234.080 7.450 234.980 ;
        RECT  1.850 234.080 3.730 234.980 ;
        RECT  1.910 0.000 32.190 4.300 ;
        LAYER metal2 ;
        POLYGON  34.100 234.980 17.650 234.980 17.650 233.800 15.210 233.800
                 15.210 234.980 11.450 234.980 11.450 233.800 9.010 233.800 9.010 234.980
                 7.730 234.980 7.730 233.800 5.290 233.800 5.290 234.980 4.010 234.980
                 4.010 233.800 1.570 233.800 1.570 234.980 0.000 234.980 0.000 0.000
                 1.590 0.000 1.590 4.620 32.510 4.620 32.510 0.000 34.100 0.000 ;
        LAYER via2 ;
        RECT  15.490 234.080 17.370 234.980 ;
        RECT  9.290 234.080 11.170 234.980 ;
        RECT  5.570 234.080 7.450 234.980 ;
        RECT  1.850 234.080 3.730 234.980 ;
        RECT  1.910 0.000 32.190 4.300 ;
        LAYER metal3 ;
        POLYGON  34.100 234.980 17.650 234.980 17.650 233.800 15.210 233.800
                 15.210 234.980 11.450 234.980 11.450 233.800 9.010 233.800 9.010 234.980
                 7.730 234.980 7.730 233.800 5.290 233.800 5.290 234.980 4.010 234.980
                 4.010 233.800 1.570 233.800 1.570 234.980 0.000 234.980 0.000 0.000
                 1.590 0.000 1.590 4.620 32.510 4.620 32.510 0.000 34.100 0.000 ;
        LAYER via3 ;
        RECT  1.910 0.000 32.190 4.300 ;
        LAYER metal4 ;
        POLYGON  34.100 234.980 0.000 234.980 0.000 0.000 1.590 0.000 1.590 4.620
                 32.510 4.620 32.510 0.000 34.100 0.000 ;
        LAYER via4 ;
        RECT  1.910 0.000 32.190 4.300 ;
        LAYER metal5 ;
        POLYGON  34.100 234.980 0.000 234.980 0.000 0.000 1.590 0.000 1.590 4.620
                 32.510 4.620 32.510 0.000 34.100 0.000 ;
        LAYER via5 ;
        RECT  1.910 0.000 32.190 4.300 ;
        LAYER metal6 ;
        POLYGON  34.100 234.980 0.000 234.980 0.000 0.000 1.310 0.000 1.310 4.900
                 32.790 4.900 32.790 0.000 34.100 0.000 ;
    END
END XMC

MACRO XMD
    CLASS PAD ;
    FOREIGN XMD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 62.620 BY 140.120 ;
    SYMMETRY x y r90 ;
    SITE iocore_d ;
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal3 ;
        RECT  39.670 138.600 41.550 139.500 ;
        LAYER metal2 ;
        RECT  39.670 138.600 41.550 139.500 ;
        LAYER metal1 ;
        RECT  39.670 138.600 41.550 139.500 ;
        END
    END O
    PIN PD
        DIRECTION INPUT ;
        PORT
        LAYER metal3 ;
        RECT  33.470 138.600 35.350 139.500 ;
        LAYER metal2 ;
        RECT  33.470 138.600 35.350 139.500 ;
        LAYER metal1 ;
        RECT  33.470 138.600 35.350 139.500 ;
        END
    END PD
    PIN SMT
        DIRECTION INPUT ;
        PORT
        LAYER metal3 ;
        RECT  23.550 138.600 25.430 139.500 ;
        LAYER metal2 ;
        RECT  23.550 138.600 25.430 139.500 ;
        LAYER metal1 ;
        RECT  23.550 138.600 25.430 139.500 ;
        END
    END SMT
    PIN PU
        DIRECTION INPUT ;
        PORT
        LAYER metal3 ;
        RECT  27.890 138.600 29.770 139.500 ;
        LAYER metal2 ;
        RECT  27.890 138.600 29.770 139.500 ;
        LAYER metal1 ;
        RECT  27.890 138.600 29.770 139.500 ;
        END
    END PU
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal6 ;
        RECT  2.850 0.000 59.770 3.000 ;
        LAYER metal5 ;
        RECT  2.850 0.000 59.770 3.000 ;
        LAYER metal4 ;
        RECT  2.850 0.000 59.770 3.000 ;
        LAYER metal3 ;
        RECT  2.850 0.000 59.770 3.000 ;
        LAYER metal2 ;
        RECT  2.850 0.000 59.770 3.000 ;
        LAYER metal1 ;
        RECT  2.850 0.000 59.770 3.000 ;
        END
    END I
    OBS
        LAYER metal1 ;
        POLYGON  62.620 139.500 41.790 139.500 41.790 138.360 39.430 138.360
                 39.430 139.500 35.590 139.500 35.590 138.360 33.230 138.360
                 33.230 139.500 30.010 139.500 30.010 138.360 27.650 138.360
                 27.650 139.500 25.670 139.500 25.670 138.360 23.310 138.360
                 23.310 139.500 0.000 139.500 0.000 0.000 2.570 0.000 2.570 3.280
                 60.050 3.280 60.050 0.000 62.620 0.000 ;
        LAYER via ;
        RECT  39.670 138.600 41.550 139.500 ;
        RECT  33.470 138.600 35.350 139.500 ;
        RECT  23.550 138.600 25.430 139.500 ;
        RECT  27.890 138.600 29.770 139.500 ;
        RECT  2.850 0.000 59.770 3.000 ;
        LAYER metal2 ;
        POLYGON  62.620 139.500 41.830 139.500 41.830 138.320 39.390 138.320
                 39.390 139.500 35.630 139.500 35.630 138.320 33.190 138.320
                 33.190 139.500 30.050 139.500 30.050 138.320 27.610 138.320
                 27.610 139.500 25.710 139.500 25.710 138.320 23.270 138.320
                 23.270 139.500 0.000 139.500 0.000 0.000 2.530 0.000 2.530 3.320
                 60.090 3.320 60.090 0.000 62.620 0.000 ;
        LAYER via2 ;
        RECT  39.670 138.600 41.550 139.500 ;
        RECT  33.470 138.600 35.350 139.500 ;
        RECT  23.550 138.600 25.430 139.500 ;
        RECT  27.890 138.600 29.770 139.500 ;
        RECT  2.850 0.000 59.770 3.000 ;
        LAYER metal3 ;
        POLYGON  62.620 139.500 41.830 139.500 41.830 138.320 39.390 138.320
                 39.390 139.500 35.630 139.500 35.630 138.320 33.190 138.320
                 33.190 139.500 30.050 139.500 30.050 138.320 27.610 138.320
                 27.610 139.500 25.710 139.500 25.710 138.320 23.270 138.320
                 23.270 139.500 0.000 139.500 0.000 0.000 2.530 0.000 2.530 3.320
                 60.090 3.320 60.090 0.000 62.620 0.000 ;
        LAYER via3 ;
        RECT  2.850 0.000 59.770 3.000 ;
        LAYER metal4 ;
        POLYGON  62.620 139.500 0.000 139.500 0.000 0.000 2.530 0.000 2.530 3.320
                 60.090 3.320 60.090 0.000 62.620 0.000 ;
        LAYER via4 ;
        RECT  2.850 0.000 59.770 3.000 ;
        LAYER metal5 ;
        POLYGON  62.620 139.500 0.000 139.500 0.000 0.000 2.530 0.000 2.530 3.320
                 60.090 3.320 60.090 0.000 62.620 0.000 ;
        LAYER via5 ;
        RECT  2.850 0.000 59.770 3.000 ;
        LAYER metal6 ;
        POLYGON  62.620 139.500 0.000 139.500 0.000 0.000 2.250 0.000 2.250 3.600
                 60.370 3.600 60.370 0.000 62.620 0.000 ;
    END
END XMD

MACRO YA2GSC
    CLASS PAD ;
    FOREIGN YA2GSC 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 34.100 BY 235.600 ;
    SYMMETRY x y r90 ;
    SITE iocore_c ;
    PIN E2
        DIRECTION INPUT ;
        PORT
        LAYER metal3 ;
        RECT  18.590 234.080 20.470 234.980 ;
        LAYER metal2 ;
        RECT  18.590 234.080 20.470 234.980 ;
        LAYER metal1 ;
        RECT  18.590 234.080 20.470 234.980 ;
        END
    END E2
    PIN E8
        DIRECTION INPUT ;
        PORT
        LAYER metal3 ;
        RECT  21.690 234.080 23.570 234.980 ;
        LAYER metal2 ;
        RECT  21.690 234.080 23.570 234.980 ;
        LAYER metal1 ;
        RECT  21.690 234.080 23.570 234.980 ;
        END
    END E8
    PIN E4
        DIRECTION INPUT ;
        PORT
        LAYER metal3 ;
        RECT  24.790 234.080 26.670 234.980 ;
        LAYER metal2 ;
        RECT  24.790 234.080 26.670 234.980 ;
        LAYER metal1 ;
        RECT  24.790 234.080 26.670 234.980 ;
        END
    END E4
    PIN SR
        DIRECTION INPUT ;
        PORT
        LAYER metal3 ;
        RECT  30.990 234.080 32.870 234.980 ;
        LAYER metal2 ;
        RECT  30.990 234.080 32.870 234.980 ;
        LAYER metal1 ;
        RECT  30.990 234.080 32.870 234.980 ;
        END
    END SR
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal3 ;
        RECT  27.890 234.080 29.770 234.980 ;
        LAYER metal2 ;
        RECT  27.890 234.080 29.770 234.980 ;
        LAYER metal1 ;
        RECT  27.890 234.080 29.770 234.980 ;
        END
    END I
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER metal3 ;
        RECT  15.490 234.080 17.370 234.980 ;
        LAYER metal2 ;
        RECT  15.490 234.080 17.370 234.980 ;
        LAYER metal1 ;
        RECT  15.490 234.080 17.370 234.980 ;
        END
    END E
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal6 ;
        RECT  1.910 0.000 32.190 4.300 ;
        LAYER metal5 ;
        RECT  1.910 0.000 32.190 4.300 ;
        LAYER metal4 ;
        RECT  1.910 0.000 32.190 4.300 ;
        LAYER metal3 ;
        RECT  1.910 0.000 32.190 4.300 ;
        LAYER metal2 ;
        RECT  1.910 0.000 32.190 4.300 ;
        LAYER metal1 ;
        RECT  1.910 0.000 32.190 4.300 ;
        END
    END O
    OBS
        LAYER metal1 ;
        POLYGON  34.100 234.980 33.110 234.980 33.110 233.840 30.750 233.840
                 30.750 234.980 30.010 234.980 30.010 233.840 27.650 233.840
                 27.650 234.980 26.910 234.980 26.910 233.840 24.550 233.840
                 24.550 234.980 23.810 234.980 23.810 233.840 21.450 233.840
                 21.450 234.980 20.710 234.980 20.710 233.840 18.350 233.840
                 18.350 234.980 17.610 234.980 17.610 233.840 15.250 233.840
                 15.250 234.980 0.000 234.980 0.000 0.000 1.630 0.000 1.630 4.580
                 32.470 4.580 32.470 0.000 34.100 0.000 ;
        LAYER via ;
        RECT  18.590 234.080 20.470 234.980 ;
        RECT  21.690 234.080 23.570 234.980 ;
        RECT  24.790 234.080 26.670 234.980 ;
        RECT  30.990 234.080 32.870 234.980 ;
        RECT  27.890 234.080 29.770 234.980 ;
        RECT  15.490 234.080 17.370 234.980 ;
        RECT  1.910 0.000 32.190 4.300 ;
        LAYER metal2 ;
        POLYGON  34.100 234.980 33.150 234.980 33.150 233.800 30.710 233.800
                 30.710 234.980 30.050 234.980 30.050 233.800 27.610 233.800
                 27.610 234.980 26.950 234.980 26.950 233.800 24.510 233.800
                 24.510 234.980 23.850 234.980 23.850 233.800 21.410 233.800
                 21.410 234.980 20.750 234.980 20.750 233.800 18.310 233.800
                 18.310 234.980 17.650 234.980 17.650 233.800 15.210 233.800
                 15.210 234.980 0.000 234.980 0.000 0.000 1.590 0.000 1.590 4.620
                 32.510 4.620 32.510 0.000 34.100 0.000 ;
        LAYER via2 ;
        RECT  18.590 234.080 20.470 234.980 ;
        RECT  21.690 234.080 23.570 234.980 ;
        RECT  24.790 234.080 26.670 234.980 ;
        RECT  30.990 234.080 32.870 234.980 ;
        RECT  27.890 234.080 29.770 234.980 ;
        RECT  15.490 234.080 17.370 234.980 ;
        RECT  1.910 0.000 32.190 4.300 ;
        LAYER metal3 ;
        POLYGON  34.100 234.980 33.150 234.980 33.150 233.800 30.710 233.800
                 30.710 234.980 30.050 234.980 30.050 233.800 27.610 233.800
                 27.610 234.980 26.950 234.980 26.950 233.800 24.510 233.800
                 24.510 234.980 23.850 234.980 23.850 233.800 21.410 233.800
                 21.410 234.980 20.750 234.980 20.750 233.800 18.310 233.800
                 18.310 234.980 17.650 234.980 17.650 233.800 15.210 233.800
                 15.210 234.980 0.000 234.980 0.000 0.000 1.590 0.000 1.590 4.620
                 32.510 4.620 32.510 0.000 34.100 0.000 ;
        LAYER via3 ;
        RECT  1.910 0.000 32.190 4.300 ;
        LAYER metal4 ;
        POLYGON  34.100 234.980 0.000 234.980 0.000 0.000 1.590 0.000 1.590 4.620
                 32.510 4.620 32.510 0.000 34.100 0.000 ;
        LAYER via4 ;
        RECT  1.910 0.000 32.190 4.300 ;
        LAYER metal5 ;
        POLYGON  34.100 234.980 0.000 234.980 0.000 0.000 1.590 0.000 1.590 4.620
                 32.510 4.620 32.510 0.000 34.100 0.000 ;
        LAYER via5 ;
        RECT  1.910 0.000 32.190 4.300 ;
        LAYER metal6 ;
        POLYGON  34.100 234.980 0.000 234.980 0.000 0.000 1.310 0.000 1.310 4.900
                 32.790 4.900 32.790 0.000 34.100 0.000 ;
    END
END YA2GSC

MACRO YA2GSD
    CLASS PAD ;
    FOREIGN YA2GSD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 62.620 BY 140.120 ;
    SYMMETRY x y r90 ;
    SITE iocore_d ;
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal3 ;
        RECT  24.170 138.600 26.050 139.500 ;
        LAYER metal2 ;
        RECT  24.170 138.600 26.050 139.500 ;
        LAYER metal1 ;
        RECT  24.170 138.600 26.050 139.500 ;
        END
    END I
    PIN E4
        DIRECTION INPUT ;
        PORT
        LAYER metal3 ;
        RECT  20.450 138.600 22.330 139.500 ;
        LAYER metal2 ;
        RECT  20.450 138.600 22.330 139.500 ;
        LAYER metal1 ;
        RECT  20.450 138.600 22.330 139.500 ;
        END
    END E4
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER metal3 ;
        RECT  33.470 138.600 35.350 139.500 ;
        LAYER metal2 ;
        RECT  33.470 138.600 35.350 139.500 ;
        LAYER metal1 ;
        RECT  33.470 138.600 35.350 139.500 ;
        END
    END E
    PIN SR
        DIRECTION INPUT ;
        PORT
        LAYER metal3 ;
        RECT  27.890 138.600 29.770 139.500 ;
        LAYER metal2 ;
        RECT  27.890 138.600 29.770 139.500 ;
        LAYER metal1 ;
        RECT  27.890 138.600 29.770 139.500 ;
        END
    END SR
    PIN E8
        DIRECTION INPUT ;
        PORT
        LAYER metal3 ;
        RECT  17.350 138.600 19.230 139.500 ;
        LAYER metal2 ;
        RECT  17.350 138.600 19.230 139.500 ;
        LAYER metal1 ;
        RECT  17.350 138.600 19.230 139.500 ;
        END
    END E8
    PIN E2
        DIRECTION INPUT ;
        PORT
        LAYER metal3 ;
        RECT  14.250 138.600 16.130 139.500 ;
        LAYER metal2 ;
        RECT  14.250 138.600 16.130 139.500 ;
        LAYER metal1 ;
        RECT  14.250 138.600 16.130 139.500 ;
        END
    END E2
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal6 ;
        RECT  2.850 0.000 59.770 3.000 ;
        LAYER metal5 ;
        RECT  2.850 0.000 59.770 3.000 ;
        LAYER metal4 ;
        RECT  2.850 0.000 59.770 3.000 ;
        LAYER metal3 ;
        RECT  2.850 0.000 59.770 3.000 ;
        LAYER metal2 ;
        RECT  2.850 0.000 59.770 3.000 ;
        LAYER metal1 ;
        RECT  2.850 0.000 59.770 3.000 ;
        END
    END O
    OBS
        LAYER metal1 ;
        POLYGON  62.620 139.500 35.590 139.500 35.590 138.360 33.230 138.360
                 33.230 139.500 30.010 139.500 30.010 138.360 27.650 138.360
                 27.650 139.500 26.290 139.500 26.290 138.360 23.930 138.360
                 23.930 139.500 22.570 139.500 22.570 138.360 20.210 138.360
                 20.210 139.500 19.470 139.500 19.470 138.360 17.110 138.360
                 17.110 139.500 16.370 139.500 16.370 138.360 14.010 138.360
                 14.010 139.500 0.000 139.500 0.000 0.000 2.570 0.000 2.570 3.280
                 60.050 3.280 60.050 0.000 62.620 0.000 ;
        LAYER via ;
        RECT  24.170 138.600 26.050 139.500 ;
        RECT  20.450 138.600 22.330 139.500 ;
        RECT  33.470 138.600 35.350 139.500 ;
        RECT  27.890 138.600 29.770 139.500 ;
        RECT  17.350 138.600 19.230 139.500 ;
        RECT  14.250 138.600 16.130 139.500 ;
        RECT  2.850 0.000 59.770 3.000 ;
        LAYER metal2 ;
        POLYGON  62.620 139.500 35.630 139.500 35.630 138.320 33.190 138.320
                 33.190 139.500 30.050 139.500 30.050 138.320 27.610 138.320
                 27.610 139.500 26.330 139.500 26.330 138.320 23.890 138.320
                 23.890 139.500 22.610 139.500 22.610 138.320 20.170 138.320
                 20.170 139.500 19.510 139.500 19.510 138.320 17.070 138.320
                 17.070 139.500 16.410 139.500 16.410 138.320 13.970 138.320
                 13.970 139.500 0.000 139.500 0.000 0.000 2.530 0.000 2.530 3.320
                 60.090 3.320 60.090 0.000 62.620 0.000 ;
        LAYER via2 ;
        RECT  24.170 138.600 26.050 139.500 ;
        RECT  20.450 138.600 22.330 139.500 ;
        RECT  33.470 138.600 35.350 139.500 ;
        RECT  27.890 138.600 29.770 139.500 ;
        RECT  17.350 138.600 19.230 139.500 ;
        RECT  14.250 138.600 16.130 139.500 ;
        RECT  2.850 0.000 59.770 3.000 ;
        LAYER metal3 ;
        POLYGON  62.620 139.500 35.630 139.500 35.630 138.320 33.190 138.320
                 33.190 139.500 30.050 139.500 30.050 138.320 27.610 138.320
                 27.610 139.500 26.330 139.500 26.330 138.320 23.890 138.320
                 23.890 139.500 22.610 139.500 22.610 138.320 20.170 138.320
                 20.170 139.500 19.510 139.500 19.510 138.320 17.070 138.320
                 17.070 139.500 16.410 139.500 16.410 138.320 13.970 138.320
                 13.970 139.500 0.000 139.500 0.000 0.000 2.530 0.000 2.530 3.320
                 60.090 3.320 60.090 0.000 62.620 0.000 ;
        LAYER via3 ;
        RECT  2.850 0.000 59.770 3.000 ;
        LAYER metal4 ;
        POLYGON  62.620 139.500 0.000 139.500 0.000 0.000 2.530 0.000 2.530 3.320
                 60.090 3.320 60.090 0.000 62.620 0.000 ;
        LAYER via4 ;
        RECT  2.850 0.000 59.770 3.000 ;
        LAYER metal5 ;
        POLYGON  62.620 139.500 0.000 139.500 0.000 0.000 2.530 0.000 2.530 3.320
                 60.090 3.320 60.090 0.000 62.620 0.000 ;
        LAYER via5 ;
        RECT  2.850 0.000 59.770 3.000 ;
        LAYER metal6 ;
        POLYGON  62.620 139.500 0.000 139.500 0.000 0.000 2.250 0.000 2.250 3.600
                 60.370 3.600 60.370 0.000 62.620 0.000 ;
    END
END YA2GSD

MACRO ZMA2GSC
    CLASS PAD ;
    FOREIGN ZMA2GSC 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 34.100 BY 235.600 ;
    SYMMETRY x y r90 ;
    SITE iocore_c ;
    PIN E2
        DIRECTION INPUT ;
        PORT
        LAYER metal3 ;
        RECT  18.590 234.080 20.470 234.980 ;
        LAYER metal2 ;
        RECT  18.590 234.080 20.470 234.980 ;
        LAYER metal1 ;
        RECT  18.590 234.080 20.470 234.980 ;
        END
    END E2
    PIN E8
        DIRECTION INPUT ;
        PORT
        LAYER metal3 ;
        RECT  21.690 234.080 23.570 234.980 ;
        LAYER metal2 ;
        RECT  21.690 234.080 23.570 234.980 ;
        LAYER metal1 ;
        RECT  21.690 234.080 23.570 234.980 ;
        END
    END E8
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal3 ;
        RECT  15.490 234.080 17.370 234.980 ;
        LAYER metal2 ;
        RECT  15.490 234.080 17.370 234.980 ;
        LAYER metal1 ;
        RECT  15.490 234.080 17.370 234.980 ;
        END
    END O
    PIN PD
        DIRECTION INPUT ;
        PORT
        LAYER metal3 ;
        RECT  9.290 234.080 11.170 234.980 ;
        LAYER metal2 ;
        RECT  9.290 234.080 11.170 234.980 ;
        LAYER metal1 ;
        RECT  9.290 234.080 11.170 234.980 ;
        END
    END PD
    PIN E4
        DIRECTION INPUT ;
        PORT
        LAYER metal3 ;
        RECT  24.790 234.080 26.670 234.980 ;
        LAYER metal2 ;
        RECT  24.790 234.080 26.670 234.980 ;
        LAYER metal1 ;
        RECT  24.790 234.080 26.670 234.980 ;
        END
    END E4
    PIN PU
        DIRECTION INPUT ;
        PORT
        LAYER metal3 ;
        RECT  5.570 234.080 7.450 234.980 ;
        LAYER metal2 ;
        RECT  5.570 234.080 7.450 234.980 ;
        LAYER metal1 ;
        RECT  5.570 234.080 7.450 234.980 ;
        END
    END PU
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER metal3 ;
        RECT  12.390 234.080 14.270 234.980 ;
        LAYER metal2 ;
        RECT  12.390 234.080 14.270 234.980 ;
        LAYER metal1 ;
        RECT  12.390 234.080 14.270 234.980 ;
        END
    END E
    PIN SR
        DIRECTION INPUT ;
        PORT
        LAYER metal3 ;
        RECT  30.990 234.080 32.870 234.980 ;
        LAYER metal2 ;
        RECT  30.990 234.080 32.870 234.980 ;
        LAYER metal1 ;
        RECT  30.990 234.080 32.870 234.980 ;
        END
    END SR
    PIN SMT
        DIRECTION INPUT ;
        PORT
        LAYER metal3 ;
        RECT  1.850 234.080 3.730 234.980 ;
        LAYER metal2 ;
        RECT  1.850 234.080 3.730 234.980 ;
        LAYER metal1 ;
        RECT  1.850 234.080 3.730 234.980 ;
        END
    END SMT
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal3 ;
        RECT  27.890 234.080 29.770 234.980 ;
        LAYER metal2 ;
        RECT  27.890 234.080 29.770 234.980 ;
        LAYER metal1 ;
        RECT  27.890 234.080 29.770 234.980 ;
        END
    END I
    PIN IO
        DIRECTION INOUT ;
        PORT
        LAYER metal6 ;
        RECT  1.910 0.000 32.190 4.300 ;
        LAYER metal5 ;
        RECT  1.910 0.000 32.190 4.300 ;
        LAYER metal4 ;
        RECT  1.910 0.000 32.190 4.300 ;
        LAYER metal3 ;
        RECT  1.910 0.000 32.190 4.300 ;
        LAYER metal2 ;
        RECT  1.910 0.000 32.190 4.300 ;
        LAYER metal1 ;
        RECT  1.910 0.000 32.190 4.300 ;
        END
    END IO
    OBS
        LAYER metal1 ;
        POLYGON  34.100 234.980 33.110 234.980 33.110 233.840 30.750 233.840
                 30.750 234.980 30.010 234.980 30.010 233.840 27.650 233.840
                 27.650 234.980 26.910 234.980 26.910 233.840 24.550 233.840
                 24.550 234.980 23.810 234.980 23.810 233.840 21.450 233.840
                 21.450 234.980 20.710 234.980 20.710 233.840 18.350 233.840
                 18.350 234.980 17.610 234.980 17.610 233.840 15.250 233.840
                 15.250 234.980 14.510 234.980 14.510 233.840 12.150 233.840
                 12.150 234.980 11.410 234.980 11.410 233.840 9.050 233.840 9.050 234.980
                 7.690 234.980 7.690 233.840 5.330 233.840 5.330 234.980 3.970 234.980
                 3.970 233.840 1.610 233.840 1.610 234.980 0.000 234.980 0.000 0.000
                 1.630 0.000 1.630 4.580 32.470 4.580 32.470 0.000 34.100 0.000 ;
        LAYER via ;
        RECT  18.590 234.080 20.470 234.980 ;
        RECT  21.690 234.080 23.570 234.980 ;
        RECT  15.490 234.080 17.370 234.980 ;
        RECT  9.290 234.080 11.170 234.980 ;
        RECT  24.790 234.080 26.670 234.980 ;
        RECT  5.570 234.080 7.450 234.980 ;
        RECT  12.390 234.080 14.270 234.980 ;
        RECT  30.990 234.080 32.870 234.980 ;
        RECT  1.850 234.080 3.730 234.980 ;
        RECT  27.890 234.080 29.770 234.980 ;
        RECT  1.910 0.000 32.190 4.300 ;
        LAYER metal2 ;
        POLYGON  34.100 234.980 33.150 234.980 33.150 233.800 30.710 233.800
                 30.710 234.980 30.050 234.980 30.050 233.800 27.610 233.800
                 27.610 234.980 26.950 234.980 26.950 233.800 24.510 233.800
                 24.510 234.980 23.850 234.980 23.850 233.800 21.410 233.800
                 21.410 234.980 20.750 234.980 20.750 233.800 18.310 233.800
                 18.310 234.980 17.650 234.980 17.650 233.800 15.210 233.800
                 15.210 234.980 14.550 234.980 14.550 233.800 12.110 233.800
                 12.110 234.980 11.450 234.980 11.450 233.800 9.010 233.800 9.010 234.980
                 7.730 234.980 7.730 233.800 5.290 233.800 5.290 234.980 4.010 234.980
                 4.010 233.800 1.570 233.800 1.570 234.980 0.000 234.980 0.000 0.000
                 1.590 0.000 1.590 4.620 32.510 4.620 32.510 0.000 34.100 0.000 ;
        LAYER via2 ;
        RECT  18.590 234.080 20.470 234.980 ;
        RECT  21.690 234.080 23.570 234.980 ;
        RECT  15.490 234.080 17.370 234.980 ;
        RECT  9.290 234.080 11.170 234.980 ;
        RECT  24.790 234.080 26.670 234.980 ;
        RECT  5.570 234.080 7.450 234.980 ;
        RECT  12.390 234.080 14.270 234.980 ;
        RECT  30.990 234.080 32.870 234.980 ;
        RECT  1.850 234.080 3.730 234.980 ;
        RECT  27.890 234.080 29.770 234.980 ;
        RECT  1.910 0.000 32.190 4.300 ;
        LAYER metal3 ;
        POLYGON  34.100 234.980 33.150 234.980 33.150 233.800 30.710 233.800
                 30.710 234.980 30.050 234.980 30.050 233.800 27.610 233.800
                 27.610 234.980 26.950 234.980 26.950 233.800 24.510 233.800
                 24.510 234.980 23.850 234.980 23.850 233.800 21.410 233.800
                 21.410 234.980 20.750 234.980 20.750 233.800 18.310 233.800
                 18.310 234.980 17.650 234.980 17.650 233.800 15.210 233.800
                 15.210 234.980 14.550 234.980 14.550 233.800 12.110 233.800
                 12.110 234.980 11.450 234.980 11.450 233.800 9.010 233.800 9.010 234.980
                 7.730 234.980 7.730 233.800 5.290 233.800 5.290 234.980 4.010 234.980
                 4.010 233.800 1.570 233.800 1.570 234.980 0.000 234.980 0.000 0.000
                 1.590 0.000 1.590 4.620 32.510 4.620 32.510 0.000 34.100 0.000 ;
        LAYER via3 ;
        RECT  1.910 0.000 32.190 4.300 ;
        LAYER metal4 ;
        POLYGON  34.100 234.980 0.000 234.980 0.000 0.000 1.590 0.000 1.590 4.620
                 32.510 4.620 32.510 0.000 34.100 0.000 ;
        LAYER via4 ;
        RECT  1.910 0.000 32.190 4.300 ;
        LAYER metal5 ;
        POLYGON  34.100 234.980 0.000 234.980 0.000 0.000 1.590 0.000 1.590 4.620
                 32.510 4.620 32.510 0.000 34.100 0.000 ;
        LAYER via5 ;
        RECT  1.910 0.000 32.190 4.300 ;
        LAYER metal6 ;
        POLYGON  34.100 234.980 0.000 234.980 0.000 0.000 1.310 0.000 1.310 4.900
                 32.790 4.900 32.790 0.000 34.100 0.000 ;
    END
END ZMA2GSC

MACRO ZMA2GSD
    CLASS PAD ;
    FOREIGN ZMA2GSD 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 62.620 BY 140.120 ;
    SYMMETRY x y r90 ;
    SITE iocore_d ;
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER metal3 ;
        RECT  32.230 138.600 34.110 139.500 ;
        LAYER metal2 ;
        RECT  32.230 138.600 34.110 139.500 ;
        LAYER metal1 ;
        RECT  32.230 138.600 34.110 139.500 ;
        END
    END I
    PIN E4
        DIRECTION INPUT ;
        PORT
        LAYER metal3 ;
        RECT  28.510 138.600 30.390 139.500 ;
        LAYER metal2 ;
        RECT  28.510 138.600 30.390 139.500 ;
        LAYER metal1 ;
        RECT  28.510 138.600 30.390 139.500 ;
        END
    END E4
    PIN O
        DIRECTION OUTPUT ;
        PORT
        LAYER metal3 ;
        RECT  17.970 138.600 19.850 139.500 ;
        LAYER metal2 ;
        RECT  17.970 138.600 19.850 139.500 ;
        LAYER metal1 ;
        RECT  17.970 138.600 19.850 139.500 ;
        END
    END O
    PIN PD
        DIRECTION INPUT ;
        PORT
        LAYER metal3 ;
        RECT  11.770 138.600 13.650 139.500 ;
        LAYER metal2 ;
        RECT  11.770 138.600 13.650 139.500 ;
        LAYER metal1 ;
        RECT  11.770 138.600 13.650 139.500 ;
        END
    END PD
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER metal3 ;
        RECT  41.530 138.600 43.410 139.500 ;
        LAYER metal2 ;
        RECT  41.530 138.600 43.410 139.500 ;
        LAYER metal1 ;
        RECT  41.530 138.600 43.410 139.500 ;
        END
    END E
    PIN SMT
        DIRECTION INPUT ;
        PORT
        LAYER metal3 ;
        RECT  1.850 138.600 3.730 139.500 ;
        LAYER metal2 ;
        RECT  1.850 138.600 3.730 139.500 ;
        LAYER metal1 ;
        RECT  1.850 138.600 3.730 139.500 ;
        END
    END SMT
    PIN PU
        DIRECTION INPUT ;
        PORT
        LAYER metal3 ;
        RECT  6.190 138.600 8.070 139.500 ;
        LAYER metal2 ;
        RECT  6.190 138.600 8.070 139.500 ;
        LAYER metal