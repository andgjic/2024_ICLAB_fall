VERSION 5.5 ;
NAMESCASESENSITIVE ON ;





LAYER metal1  
    AntennaAreaRatio 400 ;
    AntennaCumAreaRatio 400 ;
    AntennaAreaFactor 1 ;  
END metal1

LAYER metal2
    AntennaAreaRatio 400 ;
    AntennaCumAreaRatio 400 ;
    AntennaAreaFactor 1 ;  
END metal2

LAYER metal3
    AntennaAreaRatio 400 ;
    AntennaCumAreaRatio 400 ;
    AntennaAreaFactor 1 ;  
END metal3

LAYER metal4  
    AntennaAreaRatio 400 ;
    AntennaCumAreaRatio 400 ;
    AntennaAreaFactor 1 ;  
END metal4

LAYER metal5  
    AntennaAreaRatio 400 ;
    AntennaCumAreaRatio 400 ;
    AntennaAreaFactor 1 ;  
END metal5

LAYER metal6
    AntennaAreaRatio 400 ;
    AntennaCumAreaRatio 400 ;
    AntennaAreaFactor 1 ;  
END metal6


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:34:03 CST 2007
#
#**********************************************************************




MACRO AN2
  PIN I1
   AntennaPartialMetalArea                    0.201400 LAYER metal1 ;
   AntennaGateArea                            0.167400 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.274794 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.195200 LAYER metal1 ;
   AntennaGateArea                            0.169200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.615836 LAYER metal1 ; 
  END I2

  PIN O
   AntennaPartialMetalArea                    0.617600 LAYER metal1 ;
   AntennaDiffArea                            1.092700 LAYER metal1 ;
  END O

END AN2


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:34:06 CST 2007
#
#**********************************************************************




MACRO AN2B1
  PIN B1
   AntennaPartialMetalArea                    1.552000 LAYER metal1 ;
   AntennaGateArea                            0.774000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.256852 LAYER metal1 ; 
  END B1

  PIN I1
   AntennaPartialMetalArea                    0.207200 LAYER metal1 ;
   AntennaGateArea                            0.187200 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.082262 LAYER metal1 ; 
  END I1

  PIN O
   AntennaPartialMetalArea                    1.058400 LAYER metal1 ;
   AntennaDiffArea                            1.722000 LAYER metal1 ;
  END O

END AN2B1


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:34:11 CST 2007
#
#**********************************************************************




MACRO AN2B1P
  PIN B1
   AntennaPartialMetalArea                    0.227200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.972227 LAYER metal1 ; 
  END B1

  PIN I1
   AntennaPartialMetalArea                    0.203200 LAYER metal1 ;
   AntennaGateArea                            0.187200 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.361110 LAYER metal1 ; 
  END I1

  PIN O
   AntennaPartialMetalArea                    0.931200 LAYER metal1 ;
   AntennaDiffArea                            2.119600 LAYER metal1 ;
  END O

END AN2B1P


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:34:14 CST 2007
#
#**********************************************************************




MACRO AN2B1S
  PIN B1
   AntennaPartialMetalArea                    0.183200 LAYER metal1 ;
   AntennaGateArea                            0.396000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.208584 LAYER metal1 ; 
  END B1

  PIN I1
   AntennaPartialMetalArea                    0.207200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.858589 LAYER metal1 ; 
  END I1

  PIN O
   AntennaPartialMetalArea                    0.911600 LAYER metal1 ;
   AntennaDiffArea                            1.192000 LAYER metal1 ;
  END O

END AN2B1S


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:34:17 CST 2007
#
#**********************************************************************




MACRO AN2B1T
  PIN B1
   AntennaPartialMetalArea                    0.286000 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.381314 LAYER metal1 ; 
  END B1

  PIN I1
   AntennaPartialMetalArea                    0.307200 LAYER metal1 ;
   AntennaGateArea                            0.396000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.069692 LAYER metal1 ; 
  END I1

  PIN O
   AntennaPartialMetalArea                    2.904400 LAYER metal1 ;
   AntennaDiffArea                            2.865400 LAYER metal1 ;
  END O

END AN2B1T


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:34:20 CST 2007
#
#**********************************************************************




MACRO AN2P
  PIN I1
   AntennaPartialMetalArea                    0.211200 LAYER metal1 ;
   AntennaGateArea                            0.187200 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.534185 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.199200 LAYER metal1 ;
   AntennaGateArea                            0.187200 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.111107 LAYER metal1 ; 
  END I2

  PIN O
   AntennaPartialMetalArea                    0.697600 LAYER metal1 ;
   AntennaDiffArea                            1.846700 LAYER metal1 ;
  END O

END AN2P


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:34:22 CST 2007
#
#**********************************************************************




MACRO AN2S
  PIN I1
   AntennaPartialMetalArea                    0.195200 LAYER metal1 ;
   AntennaGateArea                            0.169200 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.144206 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.212800 LAYER metal1 ;
   AntennaGateArea                            0.169200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.569737 LAYER metal1 ; 
  END I2

  PIN O
   AntennaPartialMetalArea                    0.612000 LAYER metal1 ;
   AntennaDiffArea                            0.588000 LAYER metal1 ;
  END O

END AN2S


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:34:25 CST 2007
#
#**********************************************************************




MACRO AN2T
  PIN I1
   AntennaPartialMetalArea                    0.244800 LAYER metal1 ;
   AntennaGateArea                            0.396000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.261618 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.303600 LAYER metal1 ;
   AntennaGateArea                            0.396000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.061613 LAYER metal1 ; 
  END I2

  PIN O
   AntennaPartialMetalArea                    2.816400 LAYER metal1 ;
   AntennaDiffArea                            2.899000 LAYER metal1 ;
  END O

END AN2T


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:34:27 CST 2007
#
#**********************************************************************




MACRO AN3
  PIN I1
   AntennaPartialMetalArea                    0.211200 LAYER metal1 ;
   AntennaGateArea                            0.169200 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.718673 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.169200 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.250588 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.169200 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.250588 LAYER metal1 ; 
  END I3

  PIN O
   AntennaPartialMetalArea                    0.617600 LAYER metal1 ;
   AntennaDiffArea                            1.533700 LAYER metal1 ;
  END O

END AN3


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:34:30 CST 2007
#
#**********************************************************************




MACRO AN3B1
  PIN B1
   AntennaPartialMetalArea                    0.227200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.642677 LAYER metal1 ; 
  END B1

  PIN I1
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.169200 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.569738 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.169200 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.621748 LAYER metal1 ; 
  END I2

  PIN O
   AntennaPartialMetalArea                    0.617600 LAYER metal1 ;
   AntennaDiffArea                            1.533700 LAYER metal1 ;
  END O

END AN3B1


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:34:33 CST 2007
#
#**********************************************************************




MACRO AN3B1P
  PIN B1
   AntennaPartialMetalArea                    0.227200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.699497 LAYER metal1 ; 
  END B1

  PIN I1
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.169200 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.484638 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.169200 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.484638 LAYER metal1 ; 
  END I2

  PIN O
   AntennaPartialMetalArea                    0.641600 LAYER metal1 ;
   AntennaDiffArea                            1.677500 LAYER metal1 ;
  END O

END AN3B1P


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:34:35 CST 2007
#
#**********************************************************************




MACRO AN3B1S
  PIN B1
   AntennaPartialMetalArea                    0.227200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.290407 LAYER metal1 ; 
  END B1

  PIN I1
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.438127 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.460857 LAYER metal1 ; 
  END I2

  PIN O
   AntennaPartialMetalArea                    0.766000 LAYER metal1 ;
   AntennaDiffArea                            0.588000 LAYER metal1 ;
  END O

END AN3B1S


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:34:38 CST 2007
#
#**********************************************************************




MACRO AN3B1T
  PIN B1
   AntennaPartialMetalArea                    0.227200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.790407 LAYER metal1 ; 
  END B1

  PIN I1
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.270000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.637036 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.267600 LAYER metal1 ;
   AntennaGateArea                            0.270000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.637039 LAYER metal1 ; 
  END I2

  PIN O
   AntennaPartialMetalArea                    1.232400 LAYER metal1 ;
   AntennaDiffArea                            2.739000 LAYER metal1 ;
  END O

END AN3B1T


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:34:41 CST 2007
#
#**********************************************************************




MACRO AN3B2
  PIN B1
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.449497 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.211200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.654037 LAYER metal1 ; 
  END B2

  PIN I1
   AntennaPartialMetalArea                    0.350400 LAYER metal1 ;
   AntennaGateArea                            0.169200 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.718678 LAYER metal1 ; 
  END I1

  PIN O
   AntennaPartialMetalArea                    0.617600 LAYER metal1 ;
   AntennaDiffArea                            1.316500 LAYER metal1 ;
  END O

END AN3B2


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:34:44 CST 2007
#
#**********************************************************************




MACRO AN3B2P
  PIN B1
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.255047 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.211200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.654037 LAYER metal1 ; 
  END B2

  PIN I1
   AntennaPartialMetalArea                    0.252800 LAYER metal1 ;
   AntennaGateArea                            0.169200 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.718680 LAYER metal1 ; 
  END I1

  PIN O
   AntennaPartialMetalArea                    0.617600 LAYER metal1 ;
   AntennaDiffArea                            1.329000 LAYER metal1 ;
  END O

END AN3B2P


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:34:47 CST 2007
#
#**********************************************************************




MACRO AN3B2S
  PIN B1
   AntennaPartialMetalArea                    0.195200 LAYER metal1 ;
   AntennaGateArea                            0.419400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.015263 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.419400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.041013 LAYER metal1 ; 
  END B2

  PIN I1
   AntennaPartialMetalArea                    0.207200 LAYER metal1 ;
   AntennaGateArea                            0.187200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.918802 LAYER metal1 ; 
  END I1

  PIN O
   AntennaPartialMetalArea                    1.092400 LAYER metal1 ;
   AntennaDiffArea                            1.411700 LAYER metal1 ;
  END O

END AN3B2S


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:34:50 CST 2007
#
#**********************************************************************




MACRO AN3B2T
  PIN B1
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.255047 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.239200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.654039 LAYER metal1 ; 
  END B2

  PIN I1
   AntennaPartialMetalArea                    0.252800 LAYER metal1 ;
   AntennaGateArea                            0.270000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.943704 LAYER metal1 ; 
  END I1

  PIN O
   AntennaPartialMetalArea                    1.122400 LAYER metal1 ;
   AntennaDiffArea                            2.664500 LAYER metal1 ;
  END O

END AN3B2T


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:34:52 CST 2007
#
#**********************************************************************




MACRO AN3P
  PIN I1
   AntennaPartialMetalArea                    0.211200 LAYER metal1 ;
   AntennaGateArea                            0.169200 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.718673 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.169200 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.302598 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.199200 LAYER metal1 ;
   AntennaGateArea                            0.169200 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.303785 LAYER metal1 ; 
  END I3

  PIN O
   AntennaPartialMetalArea                    0.697600 LAYER metal1 ;
   AntennaDiffArea                            1.721500 LAYER metal1 ;
  END O

END AN3P


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:34:55 CST 2007
#
#**********************************************************************




MACRO AN3S
  PIN I1
   AntennaPartialMetalArea                    0.219200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.984852 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.540407 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.540407 LAYER metal1 ; 
  END I3

  PIN O
   AntennaPartialMetalArea                    0.928400 LAYER metal1 ;
   AntennaDiffArea                            0.588000 LAYER metal1 ;
  END O

END AN3S


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:34:58 CST 2007
#
#**********************************************************************




MACRO AN3T
  PIN I1
   AntennaPartialMetalArea                    0.211200 LAYER metal1 ;
   AntennaGateArea                            0.271800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.937458 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.196000 LAYER metal1 ;
   AntennaGateArea                            0.271800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.678442 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.219200 LAYER metal1 ;
   AntennaGateArea                            0.271800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.646065 LAYER metal1 ; 
  END I3

  PIN O
   AntennaPartialMetalArea                    1.218400 LAYER metal1 ;
   AntennaDiffArea                            3.223900 LAYER metal1 ;
  END O

END AN3T


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:35:02 CST 2007
#
#**********************************************************************




MACRO AN4
  PIN I1
   AntennaPartialMetalArea                    0.235600 LAYER metal1 ;
   AntennaGateArea                            0.360000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.325556 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.255200 LAYER metal1 ;
   AntennaGateArea                            0.360000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.211671 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.195200 LAYER metal1 ;
   AntennaGateArea                            0.360000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.267778 LAYER metal1 ; 
  END I3

  PIN I4
   AntennaPartialMetalArea                    0.255600 LAYER metal1 ;
   AntennaGateArea                            0.360000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.267780 LAYER metal1 ; 
  END I4

  PIN O
   AntennaPartialMetalArea                    0.846400 LAYER metal1 ;
   AntennaDiffArea                            1.657800 LAYER metal1 ;
  END O

END AN4


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:35:04 CST 2007
#
#**********************************************************************




MACRO AN4B1
  PIN B1
   AntennaPartialMetalArea                    1.427600 LAYER metal1 ;
   AntennaGateArea                            0.879600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.070460 LAYER metal1 ; 
  END B1

  PIN I1
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.439800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.947702 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.298400 LAYER metal1 ;
   AntennaGateArea                            0.438600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.010483 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.195200 LAYER metal1 ;
   AntennaGateArea                            0.438600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.301418 LAYER metal1 ; 
  END I3

  PIN O
   AntennaPartialMetalArea                    0.732400 LAYER metal1 ;
   AntennaDiffArea                            1.927000 LAYER metal1 ;
  END O

END AN4B1


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:35:07 CST 2007
#
#**********************************************************************




MACRO AN4B1P
  PIN B1
   AntennaPartialMetalArea                    1.127200 LAYER metal1 ;
   AntennaGateArea                            1.749600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.087598 LAYER metal1 ; 
  END B1

  PIN I1
   AntennaPartialMetalArea                    0.215200 LAYER metal1 ;
   AntennaGateArea                            0.542400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.707595 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.249200 LAYER metal1 ;
   AntennaGateArea                            0.537600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.664808 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.195200 LAYER metal1 ;
   AntennaGateArea                            0.547200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.998905 LAYER metal1 ; 
  END I3

  PIN O
   AntennaPartialMetalArea                    2.469600 LAYER metal1 ;
   AntennaDiffArea                            3.692400 LAYER metal1 ;
  END O

END AN4B1P


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:35:10 CST 2007
#
#**********************************************************************




MACRO AN4B1S
  PIN B1
   AntennaPartialMetalArea                    0.221600 LAYER metal1 ;
   AntennaGateArea                            0.342000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.859647 LAYER metal1 ; 
  END B1

  PIN I1
   AntennaPartialMetalArea                    0.187200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.119952 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.228000 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.483586 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.219200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.758842 LAYER metal1 ; 
  END I3

  PIN O
   AntennaPartialMetalArea                    1.372800 LAYER metal1 ;
   AntennaDiffArea                            1.211000 LAYER metal1 ;
  END O

END AN4B1S


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:35:13 CST 2007
#
#**********************************************************************




MACRO AN4B1T
  PIN B1
   AntennaPartialMetalArea                    2.572000 LAYER metal1 ;
   AntennaGateArea                            2.649600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.078347 LAYER metal1 ; 
  END B1

  PIN I1
   AntennaPartialMetalArea                    0.187200 LAYER metal1 ;
   AntennaGateArea                            0.527400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.660601 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.223200 LAYER metal1 ;
   AntennaGateArea                            0.527400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.660602 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.219200 LAYER metal1 ;
   AntennaGateArea                            0.527400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.660596 LAYER metal1 ; 
  END I3

  PIN O
   AntennaPartialMetalArea                    3.200000 LAYER metal1 ;
   AntennaDiffArea                            5.811600 LAYER metal1 ;
  END O

END AN4B1T


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:35:16 CST 2007
#
#**********************************************************************




MACRO AN4P
  PIN I1
   AntennaPartialMetalArea                    0.227200 LAYER metal1 ;
   AntennaGateArea                            0.513600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.873052 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.219200 LAYER metal1 ;
   AntennaGateArea                            0.504000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.814679 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.187200 LAYER metal1 ;
   AntennaGateArea                            0.500400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.750199 LAYER metal1 ; 
  END I3

  PIN I4
   AntennaPartialMetalArea                    0.223200 LAYER metal1 ;
   AntennaGateArea                            0.500400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.785367 LAYER metal1 ; 
  END I4

  PIN O
   AntennaPartialMetalArea                    2.971600 LAYER metal1 ;
   AntennaDiffArea                            3.747950 LAYER metal1 ;
  END O

END AN4P


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:35:18 CST 2007
#
#**********************************************************************




MACRO AN4S
  PIN I1
   AntennaPartialMetalArea                    0.199200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.450754 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.237200 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.108585 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.184800 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          4.040403 LAYER metal1 ; 
  END I3

  PIN I4
   AntennaPartialMetalArea                    0.202400 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.753792 LAYER metal1 ; 
  END I4

  PIN O
   AntennaPartialMetalArea                    1.102800 LAYER metal1 ;
   AntennaDiffArea                            0.956000 LAYER metal1 ;
  END O

END AN4S


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:35:21 CST 2007
#
#**********************************************************************




MACRO AN4T
  PIN I1
   AntennaPartialMetalArea                    0.227200 LAYER metal1 ;
   AntennaGateArea                            0.513600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.873052 LAYER metal1 ; 
  END I1

  PIN I2
   AntennaPartialMetalArea                    0.219200 LAYER metal1 ;
   AntennaGateArea                            0.504000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.814679 LAYER metal1 ; 
  END I2

  PIN I3
   AntennaPartialMetalArea                    0.187200 LAYER metal1 ;
   AntennaGateArea                            0.500400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.750199 LAYER metal1 ; 
  END I3

  PIN I4
   AntennaPartialMetalArea                    0.223200 LAYER metal1 ;
   AntennaGateArea                            0.500400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.785367 LAYER metal1 ; 
  END I4

  PIN O
   AntennaPartialMetalArea                    3.324800 LAYER metal1 ;
   AntennaDiffArea                            5.811600 LAYER metal1 ;
  END O

END AN4T


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:35:24 CST 2007
#
#**********************************************************************




MACRO ANTENNA
  PIN A
   AntennaPartialMetalArea                    0.396000 LAYER metal1 ;
   AntennaDiffArea                            0.360000 LAYER metal1 ;
  END A

END ANTENNA


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:35:27 CST 2007
#
#**********************************************************************




MACRO AO112
  PIN A1
   AntennaPartialMetalArea                    0.198000 LAYER metal1 ;
   AntennaGateArea                            0.345600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.667823 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.202400 LAYER metal1 ;
   AntennaGateArea                            0.345600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.591432 LAYER metal1 ; 
  END B1

  PIN C1
   AntennaPartialMetalArea                    0.202000 LAYER metal1 ;
   AntennaGateArea                            0.385200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.286087 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.182000 LAYER metal1 ;
   AntennaGateArea                            0.385200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.303218 LAYER metal1 ; 
  END C2

  PIN O
   AntennaPartialMetalArea                    0.553200 LAYER metal1 ;
   AntennaDiffArea                            1.363750 LAYER metal1 ;
  END O

END AO112


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:35:29 CST 2007
#
#**********************************************************************




MACRO AO112P
  PIN A1
   AntennaPartialMetalArea                    0.276400 LAYER metal1 ;
   AntennaGateArea                            0.437400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.017834 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.304400 LAYER metal1 ;
   AntennaGateArea                            0.378000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.608469 LAYER metal1 ; 
  END B1

  PIN C1
   AntennaPartialMetalArea                    0.263200 LAYER metal1 ;
   AntennaGateArea                            0.473400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.735952 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.295200 LAYER metal1 ;
   AntennaGateArea                            0.473400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.758766 LAYER metal1 ; 
  END C2

  PIN O
   AntennaPartialMetalArea                    0.902000 LAYER metal1 ;
   AntennaDiffArea                            1.690200 LAYER metal1 ;
  END O

END AO112P


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:35:32 CST 2007
#
#**********************************************************************




MACRO AO112S
  PIN A1
   AntennaPartialMetalArea                    0.222000 LAYER metal1 ;
   AntennaGateArea                            0.241200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.774462 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.186000 LAYER metal1 ;
   AntennaGateArea                            0.241200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.847426 LAYER metal1 ; 
  END B1

  PIN C1
   AntennaPartialMetalArea                    0.182000 LAYER metal1 ;
   AntennaGateArea                            0.241200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.362359 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.182000 LAYER metal1 ;
   AntennaGateArea                            0.241200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.481759 LAYER metal1 ; 
  END C2

  PIN O
   AntennaPartialMetalArea                    0.853600 LAYER metal1 ;
   AntennaDiffArea                            0.661000 LAYER metal1 ;
  END O

END AO112S


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:35:35 CST 2007
#
#**********************************************************************




MACRO AO112T
  PIN A1
   AntennaPartialMetalArea                    0.276400 LAYER metal1 ;
   AntennaGateArea                            0.437400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.017834 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.307200 LAYER metal1 ;
   AntennaGateArea                            0.378000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.526982 LAYER metal1 ; 
  END B1

  PIN C1
   AntennaPartialMetalArea                    0.291200 LAYER metal1 ;
   AntennaGateArea                            0.473400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.735955 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.267200 LAYER metal1 ;
   AntennaGateArea                            0.473400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.791722 LAYER metal1 ; 
  END C2

  PIN O
   AntennaPartialMetalArea                    1.252400 LAYER metal1 ;
   AntennaDiffArea                            3.223900 LAYER metal1 ;
  END O

END AO112T


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:35:38 CST 2007
#
#**********************************************************************




MACRO AO12
  PIN A1
   AntennaPartialMetalArea                    0.225200 LAYER metal1 ;
   AntennaGateArea                            0.241200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.377285 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.261200 LAYER metal1 ;
   AntennaGateArea                            0.270000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.065923 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.245600 LAYER metal1 ;
   AntennaGateArea                            0.270000 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.505930 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    0.799600 LAYER metal1 ;
   AntennaDiffArea                            1.556300 LAYER metal1 ;
  END O

END AO12


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:35:41 CST 2007
#
#**********************************************************************




MACRO AO12P
  PIN A1
   AntennaPartialMetalArea                    0.225200 LAYER metal1 ;
   AntennaGateArea                            0.324000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.503088 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.261200 LAYER metal1 ;
   AntennaGateArea                            0.360000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.299444 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.195200 LAYER metal1 ;
   AntennaGateArea                            0.360000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.629448 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    0.682800 LAYER metal1 ;
   AntennaDiffArea                            1.672400 LAYER metal1 ;
  END O

END AO12P


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:35:44 CST 2007
#
#**********************************************************************




MACRO AO12S
  PIN A1
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.198000 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.095959 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.223600 LAYER metal1 ;
   AntennaGateArea                            0.198000 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.358587 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.209200 LAYER metal1 ;
   AntennaGateArea                            0.198000 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.780804 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    0.852800 LAYER metal1 ;
   AntennaDiffArea                            0.588000 LAYER metal1 ;
  END O

END AO12S


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:35:47 CST 2007
#
#**********************************************************************




MACRO AO12T
  PIN A1
   AntennaPartialMetalArea                    0.225200 LAYER metal1 ;
   AntennaGateArea                            0.509400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.683941 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.261200 LAYER metal1 ;
   AntennaGateArea                            0.563400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.680866 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.251200 LAYER metal1 ;
   AntennaGateArea                            0.563400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.790206 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    1.293200 LAYER metal1 ;
   AntennaDiffArea                            2.973700 LAYER metal1 ;
  END O

END AO12T


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:35:49 CST 2007
#
#**********************************************************************




MACRO AO13
  PIN A1
   AntennaPartialMetalArea                    0.190400 LAYER metal1 ;
   AntennaGateArea                            0.295200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.795054 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.197200 LAYER metal1 ;
   AntennaGateArea                            0.396000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.052530 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.396000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.052525 LAYER metal1 ; 
  END B2

  PIN B3
   AntennaPartialMetalArea                    0.252000 LAYER metal1 ;
   AntennaGateArea                            0.396000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.374746 LAYER metal1 ; 
  END B3

  PIN O
   AntennaPartialMetalArea                    0.718400 LAYER metal1 ;
   AntennaDiffArea                            1.636950 LAYER metal1 ;
  END O

END AO13


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:35:52 CST 2007
#
#**********************************************************************




MACRO AO13P
  PIN A1
   AntennaPartialMetalArea                    0.225200 LAYER metal1 ;
   AntennaGateArea                            0.455400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.021520 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.234600 LAYER metal1 ;
   AntennaGateArea                            0.563400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.618390 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.191200 LAYER metal1 ;
   AntennaGateArea                            0.563400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.618389 LAYER metal1 ; 
  END B2

  PIN B3
   AntennaPartialMetalArea                    0.252000 LAYER metal1 ;
   AntennaGateArea                            0.563400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.790206 LAYER metal1 ; 
  END B3

  PIN O
   AntennaPartialMetalArea                    0.900800 LAYER metal1 ;
   AntennaDiffArea                            1.739600 LAYER metal1 ;
  END O

END AO13P


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:35:55 CST 2007
#
#**********************************************************************




MACRO AO13S
  PIN A1
   AntennaPartialMetalArea                    0.185600 LAYER metal1 ;
   AntennaGateArea                            0.158400 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.233583 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.209200 LAYER metal1 ;
   AntennaGateArea                            0.187200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.830129 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.202400 LAYER metal1 ;
   AntennaGateArea                            0.187200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.736113 LAYER metal1 ; 
  END B2

  PIN B3
   AntennaPartialMetalArea                    0.186000 LAYER metal1 ;
   AntennaGateArea                            0.187200 LAYER metal1 ;
   AntennaMaxAreaCAR                          3.300210 LAYER metal1 ; 
  END B3

  PIN O
   AntennaPartialMetalArea                    0.960400 LAYER metal1 ;
   AntennaDiffArea                            0.614200 LAYER metal1 ;
  END O

END AO13S


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:35:57 CST 2007
#
#**********************************************************************




MACRO AO13T
  PIN A1
   AntennaPartialMetalArea                    0.281200 LAYER metal1 ;
   AntennaGateArea                            0.455400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.021521 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.302600 LAYER metal1 ;
   AntennaGateArea                            0.563400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.618384 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.249200 LAYER metal1 ;
   AntennaGateArea                            0.563400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.618385 LAYER metal1 ; 
  END B2

  PIN B3
   AntennaPartialMetalArea                    0.279000 LAYER metal1 ;
   AntennaGateArea                            0.563400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.790202 LAYER metal1 ; 
  END B3

  PIN O
   AntennaPartialMetalArea                    1.198400 LAYER metal1 ;
   AntennaDiffArea                            3.063950 LAYER metal1 ;
  END O

END AO13T


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:36:00 CST 2007
#
#**********************************************************************




MACRO AO22
  PIN A1
   AntennaPartialMetalArea                    0.182000 LAYER metal1 ;
   AntennaGateArea                            0.327000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.533335 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.190000 LAYER metal1 ;
   AntennaGateArea                            0.327000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.555350 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.182000 LAYER metal1 ;
   AntennaGateArea                            0.322200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.533833 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.209600 LAYER metal1 ;
   AntennaGateArea                            0.322200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.902542 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    0.500000 LAYER metal1 ;
   AntennaDiffArea                            1.280450 LAYER metal1 ;
  END O

END AO22


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:36:03 CST 2007
#
#**********************************************************************




MACRO AO222
  PIN A1
   AntennaPartialMetalArea                    0.251600 LAYER metal1 ;
   AntennaGateArea                            0.384600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.188244 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.183200 LAYER metal1 ;
   AntennaGateArea                            0.384600 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.149251 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.272000 LAYER metal1 ;
   AntennaGateArea                            0.386400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.178056 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.196000 LAYER metal1 ;
   AntennaGateArea                            0.382800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.281083 LAYER metal1 ; 
  END B2

  PIN C1
   AntennaPartialMetalArea                    0.214000 LAYER metal1 ;
   AntennaGateArea                            0.390000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.437952 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.240000 LAYER metal1 ;
   AntennaGateArea                            0.390000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.133335 LAYER metal1 ; 
  END C2

  PIN O
   AntennaPartialMetalArea                    0.550400 LAYER metal1 ;
   AntennaDiffArea                            1.254950 LAYER metal1 ;
  END O

END AO222


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:36:06 CST 2007
#
#**********************************************************************




MACRO AO222P
  PIN A1
   AntennaPartialMetalArea                    0.199600 LAYER metal1 ;
   AntennaGateArea                            0.463800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.914192 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.196000 LAYER metal1 ;
   AntennaGateArea                            0.455400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.022619 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.212000 LAYER metal1 ;
   AntennaGateArea                            0.459600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.981289 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.196000 LAYER metal1 ;
   AntennaGateArea                            0.453600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.934741 LAYER metal1 ; 
  END B2

  PIN C1
   AntennaPartialMetalArea                    0.214000 LAYER metal1 ;
   AntennaGateArea                            0.458400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.184119 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.244000 LAYER metal1 ;
   AntennaGateArea                            0.458400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.924954 LAYER metal1 ; 
  END C2

  PIN O
   AntennaPartialMetalArea                    0.854000 LAYER metal1 ;
   AntennaDiffArea                            1.606500 LAYER metal1 ;
  END O

END AO222P


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:36:09 CST 2007
#
#**********************************************************************




MACRO AO222S
  PIN A1
   AntennaPartialMetalArea                    0.191600 LAYER metal1 ;
   AntennaGateArea                            0.309000 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.680905 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.183200 LAYER metal1 ;
   AntennaGateArea                            0.295200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.765584 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.196000 LAYER metal1 ;
   AntennaGateArea                            0.307200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.690759 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.196000 LAYER metal1 ;
   AntennaGateArea                            0.295200 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.759483 LAYER metal1 ; 
  END B2

  PIN C1
   AntennaPartialMetalArea                    0.214000 LAYER metal1 ;
   AntennaGateArea                            0.295200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.161928 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.240000 LAYER metal1 ;
   AntennaGateArea                            0.304800 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.704068 LAYER metal1 ; 
  END C2

  PIN O
   AntennaPartialMetalArea                    0.796800 LAYER metal1 ;
   AntennaDiffArea                            0.603000 LAYER metal1 ;
  END O

END AO222S


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:36:12 CST 2007
#
#**********************************************************************




MACRO AO222T
  PIN A1
   AntennaPartialMetalArea                    0.227600 LAYER metal1 ;
   AntennaGateArea                            0.517800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.730008 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.248400 LAYER metal1 ;
   AntennaGateArea                            0.509400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.789167 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.248400 LAYER metal1 ;
   AntennaGateArea                            0.519000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.764937 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.196000 LAYER metal1 ;
   AntennaGateArea                            0.516600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.716226 LAYER metal1 ; 
  END B2

  PIN C1
   AntennaPartialMetalArea                    0.214000 LAYER metal1 ;
   AntennaGateArea                            0.517800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.943993 LAYER metal1 ; 
  END C1

  PIN C2
   AntennaPartialMetalArea                    0.280400 LAYER metal1 ;
   AntennaGateArea                            0.517800 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.714558 LAYER metal1 ; 
  END C2

  PIN O
   AntennaPartialMetalArea                    1.246000 LAYER metal1 ;
   AntennaDiffArea                            2.747450 LAYER metal1 ;
  END O

END AO222T


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:36:15 CST 2007
#
#**********************************************************************




MACRO AO22P
  PIN A1
   AntennaPartialMetalArea                    0.217600 LAYER metal1 ;
   AntennaGateArea                            0.489000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.797140 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.177600 LAYER metal1 ;
   AntennaGateArea                            0.489000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.833130 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.217600 LAYER metal1 ;
   AntennaGateArea                            0.494400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.784791 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.206400 LAYER metal1 ;
   AntennaGateArea                            0.494400 LAYER metal1 ;
   AntennaMaxAreaCAR                          1.042884 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    0.640000 LAYER metal1 ;
   AntennaDiffArea                            1.799850 LAYER metal1 ;
  END O

END AO22P


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:36:19 CST 2007
#
#**********************************************************************




MACRO AO22S
  PIN A1
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.241200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.198178 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.204400 LAYER metal1 ;
   AntennaGateArea                            0.241200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.198180 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            0.241200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.522388 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.195200 LAYER metal1 ;
   AntennaGateArea                            0.241200 LAYER metal1 ;
   AntennaMaxAreaCAR                          2.923713 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    0.799600 LAYER metal1 ;
   AntennaDiffArea                            0.588000 LAYER metal1 ;
  END O

END AO22S


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:36:21 CST 2007
#
#**********************************************************************




MACRO AO22T
  PIN A1
   AntennaPartialMetalArea                    0.233600 LAYER metal1 ;
   AntennaGateArea                            0.561000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.624241 LAYER metal1 ; 
  END A1

  PIN A2
   AntennaPartialMetalArea                    0.193600 LAYER metal1 ;
   AntennaGateArea                            0.561000 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.655612 LAYER metal1 ; 
  END A2

  PIN B1
   AntennaPartialMetalArea                    0.217600 LAYER metal1 ;
   AntennaGateArea                            0.567600 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.613812 LAYER metal1 ; 
  END B1

  PIN B2
   AntennaPartialMetalArea                    0.224400 LAYER metal1 ;
   AntennaGateArea                            0.566400 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.832624 LAYER metal1 ; 
  END B2

  PIN O
   AntennaPartialMetalArea                    1.205600 LAYER metal1 ;
   AntennaDiffArea                            2.998400 LAYER metal1 ;
  END O

END AO22T


#**********************************************************************
#
# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
#
# Generated by Calibre Antenna verification/extraction utility antEx
#
# Gen-Date: Tue Nov  6 17:36:24 CST 2007
#
#**********************************************************************




MACRO AOI112H
  PIN A1
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            1.528200 LAYER metal1 ;
   AntennaMaxAreaCAR                          0.770318 LAYER metal1 ; 
  END A1

  PIN B1
   AntennaPartialMetalArea                    0.179200 LAYER metal1 ;
   AntennaGateArea                            1.528200 LAYER metal1 ;
   AntennaMaxAreaCAR