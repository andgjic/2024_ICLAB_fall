# 
#              Synchronous Dual Port SRAM Compiler 
# 
#                    UMC 0.18um Generic Logic Process 
#    __________________________________________________________________________
# 
# 
#      (C) Copyright 2002-2009 Faraday Technology Corp. All Rights Reserved.
#    
#    This source code is an unpublished work belongs to Faraday Technology
#    Corp.  It is considered a trade secret and is not to be divulged or
#    used by parties who have not received written authorization from
#    Faraday Technology Corp.
#    
#    Faraday's home page can be found at:
#    http://www.faraday-tech.com/
#   
#       Module Name      : DPSRAM_32_256
#       Words            : 256
#       Bits             : 32
#       Byte-Write       : 1
#       Aspect Ratio     : 1
#       Output Loading   : 0.05  (pf)
#       Data Slew        : 0.02  (ns)
#       CK Slew          : 0.02  (ns)
#       Power Ring Width : 2  (um)
# 
# -----------------------------------------------------------------------------
# 
#       Library          : FSA0M_A
#       Memaker          : 200901.2.1
#       Date             : 2024/10/28 14:00:14
# 
# -----------------------------------------------------------------------------


NAMESCASESENSITIVE ON ;
MACRO DPSRAM_32_256
CLASS BLOCK ;
FOREIGN DPSRAM_32_256 0.000 0.000 ;
ORIGIN 0.000 0.000 ;
SIZE 972.780 BY 252.560 ;
SYMMETRY x y r90 ;
SITE core ;
PIN GND
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
 PORT
  LAYER ME5 ;
  RECT 971.660 207.540 972.780 210.780 ;
  LAYER ME4 ;
  RECT 971.660 207.540 972.780 210.780 ;
  LAYER ME3 ;
  RECT 971.660 207.540 972.780 210.780 ;
  LAYER ME2 ;
  RECT 971.660 207.540 972.780 210.780 ;
  LAYER ME1 ;
  RECT 971.660 207.540 972.780 210.780 ;
 END
 PORT
  LAYER ME5 ;
  RECT 971.660 199.700 972.780 202.940 ;
  LAYER ME4 ;
  RECT 971.660 199.700 972.780 202.940 ;
  LAYER ME3 ;
  RECT 971.660 199.700 972.780 202.940 ;
  LAYER ME2 ;
  RECT 971.660 199.700 972.780 202.940 ;
  LAYER ME1 ;
  RECT 971.660 199.700 972.780 202.940 ;
 END
 PORT
  LAYER ME5 ;
  RECT 971.660 191.860 972.780 195.100 ;
  LAYER ME4 ;
  RECT 971.660 191.860 972.780 195.100 ;
  LAYER ME3 ;
  RECT 971.660 191.860 972.780 195.100 ;
  LAYER ME2 ;
  RECT 971.660 191.860 972.780 195.100 ;
  LAYER ME1 ;
  RECT 971.660 191.860 972.780 195.100 ;
 END
 PORT
  LAYER ME5 ;
  RECT 971.660 184.020 972.780 187.260 ;
  LAYER ME4 ;
  RECT 971.660 184.020 972.780 187.260 ;
  LAYER ME3 ;
  RECT 971.660 184.020 972.780 187.260 ;
  LAYER ME2 ;
  RECT 971.660 184.020 972.780 187.260 ;
  LAYER ME1 ;
  RECT 971.660 184.020 972.780 187.260 ;
 END
 PORT
  LAYER ME5 ;
  RECT 971.660 176.180 972.780 179.420 ;
  LAYER ME4 ;
  RECT 971.660 176.180 972.780 179.420 ;
  LAYER ME3 ;
  RECT 971.660 176.180 972.780 179.420 ;
  LAYER ME2 ;
  RECT 971.660 176.180 972.780 179.420 ;
  LAYER ME1 ;
  RECT 971.660 176.180 972.780 179.420 ;
 END
 PORT
  LAYER ME5 ;
  RECT 971.660 168.340 972.780 171.580 ;
  LAYER ME4 ;
  RECT 971.660 168.340 972.780 171.580 ;
  LAYER ME3 ;
  RECT 971.660 168.340 972.780 171.580 ;
  LAYER ME2 ;
  RECT 971.660 168.340 972.780 171.580 ;
  LAYER ME1 ;
  RECT 971.660 168.340 972.780 171.580 ;
 END
 PORT
  LAYER ME5 ;
  RECT 971.660 129.140 972.780 132.380 ;
  LAYER ME4 ;
  RECT 971.660 129.140 972.780 132.380 ;
  LAYER ME3 ;
  RECT 971.660 129.140 972.780 132.380 ;
  LAYER ME2 ;
  RECT 971.660 129.140 972.780 132.380 ;
  LAYER ME1 ;
  RECT 971.660 129.140 972.780 132.380 ;
 END
 PORT
  LAYER ME5 ;
  RECT 971.660 121.300 972.780 124.540 ;
  LAYER ME4 ;
  RECT 971.660 121.300 972.780 124.540 ;
  LAYER ME3 ;
  RECT 971.660 121.300 972.780 124.540 ;
  LAYER ME2 ;
  RECT 971.660 121.300 972.780 124.540 ;
  LAYER ME1 ;
  RECT 971.660 121.300 972.780 124.540 ;
 END
 PORT
  LAYER ME5 ;
  RECT 971.660 113.460 972.780 116.700 ;
  LAYER ME4 ;
  RECT 971.660 113.460 972.780 116.700 ;
  LAYER ME3 ;
  RECT 971.660 113.460 972.780 116.700 ;
  LAYER ME2 ;
  RECT 971.660 113.460 972.780 116.700 ;
  LAYER ME1 ;
  RECT 971.660 113.460 972.780 116.700 ;
 END
 PORT
  LAYER ME5 ;
  RECT 971.660 105.620 972.780 108.860 ;
  LAYER ME4 ;
  RECT 971.660 105.620 972.780 108.860 ;
  LAYER ME3 ;
  RECT 971.660 105.620 972.780 108.860 ;
  LAYER ME2 ;
  RECT 971.660 105.620 972.780 108.860 ;
  LAYER ME1 ;
  RECT 971.660 105.620 972.780 108.860 ;
 END
 PORT
  LAYER ME5 ;
  RECT 971.660 97.780 972.780 101.020 ;
  LAYER ME4 ;
  RECT 971.660 97.780 972.780 101.020 ;
  LAYER ME3 ;
  RECT 971.660 97.780 972.780 101.020 ;
  LAYER ME2 ;
  RECT 971.660 97.780 972.780 101.020 ;
  LAYER ME1 ;
  RECT 971.660 97.780 972.780 101.020 ;
 END
 PORT
  LAYER ME5 ;
  RECT 971.660 89.940 972.780 93.180 ;
  LAYER ME4 ;
  RECT 971.660 89.940 972.780 93.180 ;
  LAYER ME3 ;
  RECT 971.660 89.940 972.780 93.180 ;
  LAYER ME2 ;
  RECT 971.660 89.940 972.780 93.180 ;
  LAYER ME1 ;
  RECT 971.660 89.940 972.780 93.180 ;
 END
 PORT
  LAYER ME5 ;
  RECT 971.660 50.740 972.780 53.980 ;
  LAYER ME4 ;
  RECT 971.660 50.740 972.780 53.980 ;
  LAYER ME3 ;
  RECT 971.660 50.740 972.780 53.980 ;
  LAYER ME2 ;
  RECT 971.660 50.740 972.780 53.980 ;
  LAYER ME1 ;
  RECT 971.660 50.740 972.780 53.980 ;
 END
 PORT
  LAYER ME5 ;
  RECT 971.660 42.900 972.780 46.140 ;
  LAYER ME4 ;
  RECT 971.660 42.900 972.780 46.140 ;
  LAYER ME3 ;
  RECT 971.660 42.900 972.780 46.140 ;
  LAYER ME2 ;
  RECT 971.660 42.900 972.780 46.140 ;
  LAYER ME1 ;
  RECT 971.660 42.900 972.780 46.140 ;
 END
 PORT
  LAYER ME5 ;
  RECT 971.660 35.060 972.780 38.300 ;
  LAYER ME4 ;
  RECT 971.660 35.060 972.780 38.300 ;
  LAYER ME3 ;
  RECT 971.660 35.060 972.780 38.300 ;
  LAYER ME2 ;
  RECT 971.660 35.060 972.780 38.300 ;
  LAYER ME1 ;
  RECT 971.660 35.060 972.780 38.300 ;
 END
 PORT
  LAYER ME5 ;
  RECT 971.660 27.220 972.780 30.460 ;
  LAYER ME4 ;
  RECT 971.660 27.220 972.780 30.460 ;
  LAYER ME3 ;
  RECT 971.660 27.220 972.780 30.460 ;
  LAYER ME2 ;
  RECT 971.660 27.220 972.780 30.460 ;
  LAYER ME1 ;
  RECT 971.660 27.220 972.780 30.460 ;
 END
 PORT
  LAYER ME5 ;
  RECT 971.660 19.380 972.780 22.620 ;
  LAYER ME4 ;
  RECT 971.660 19.380 972.780 22.620 ;
  LAYER ME3 ;
  RECT 971.660 19.380 972.780 22.620 ;
  LAYER ME2 ;
  RECT 971.660 19.380 972.780 22.620 ;
  LAYER ME1 ;
  RECT 971.660 19.380 972.780 22.620 ;
 END
 PORT
  LAYER ME5 ;
  RECT 971.660 11.540 972.780 14.780 ;
  LAYER ME4 ;
  RECT 971.660 11.540 972.780 14.780 ;
  LAYER ME3 ;
  RECT 971.660 11.540 972.780 14.780 ;
  LAYER ME2 ;
  RECT 971.660 11.540 972.780 14.780 ;
  LAYER ME1 ;
  RECT 971.660 11.540 972.780 14.780 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 207.540 1.120 210.780 ;
  LAYER ME4 ;
  RECT 0.000 207.540 1.120 210.780 ;
  LAYER ME3 ;
  RECT 0.000 207.540 1.120 210.780 ;
  LAYER ME2 ;
  RECT 0.000 207.540 1.120 210.780 ;
  LAYER ME1 ;
  RECT 0.000 207.540 1.120 210.780 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 199.700 1.120 202.940 ;
  LAYER ME4 ;
  RECT 0.000 199.700 1.120 202.940 ;
  LAYER ME3 ;
  RECT 0.000 199.700 1.120 202.940 ;
  LAYER ME2 ;
  RECT 0.000 199.700 1.120 202.940 ;
  LAYER ME1 ;
  RECT 0.000 199.700 1.120 202.940 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 191.860 1.120 195.100 ;
  LAYER ME4 ;
  RECT 0.000 191.860 1.120 195.100 ;
  LAYER ME3 ;
  RECT 0.000 191.860 1.120 195.100 ;
  LAYER ME2 ;
  RECT 0.000 191.860 1.120 195.100 ;
  LAYER ME1 ;
  RECT 0.000 191.860 1.120 195.100 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 184.020 1.120 187.260 ;
  LAYER ME4 ;
  RECT 0.000 184.020 1.120 187.260 ;
  LAYER ME3 ;
  RECT 0.000 184.020 1.120 187.260 ;
  LAYER ME2 ;
  RECT 0.000 184.020 1.120 187.260 ;
  LAYER ME1 ;
  RECT 0.000 184.020 1.120 187.260 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 176.180 1.120 179.420 ;
  LAYER ME4 ;
  RECT 0.000 176.180 1.120 179.420 ;
  LAYER ME3 ;
  RECT 0.000 176.180 1.120 179.420 ;
  LAYER ME2 ;
  RECT 0.000 176.180 1.120 179.420 ;
  LAYER ME1 ;
  RECT 0.000 176.180 1.120 179.420 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 168.340 1.120 171.580 ;
  LAYER ME4 ;
  RECT 0.000 168.340 1.120 171.580 ;
  LAYER ME3 ;
  RECT 0.000 168.340 1.120 171.580 ;
  LAYER ME2 ;
  RECT 0.000 168.340 1.120 171.580 ;
  LAYER ME1 ;
  RECT 0.000 168.340 1.120 171.580 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 129.140 1.120 132.380 ;
  LAYER ME4 ;
  RECT 0.000 129.140 1.120 132.380 ;
  LAYER ME3 ;
  RECT 0.000 129.140 1.120 132.380 ;
  LAYER ME2 ;
  RECT 0.000 129.140 1.120 132.380 ;
  LAYER ME1 ;
  RECT 0.000 129.140 1.120 132.380 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 121.300 1.120 124.540 ;
  LAYER ME4 ;
  RECT 0.000 121.300 1.120 124.540 ;
  LAYER ME3 ;
  RECT 0.000 121.300 1.120 124.540 ;
  LAYER ME2 ;
  RECT 0.000 121.300 1.120 124.540 ;
  LAYER ME1 ;
  RECT 0.000 121.300 1.120 124.540 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 113.460 1.120 116.700 ;
  LAYER ME4 ;
  RECT 0.000 113.460 1.120 116.700 ;
  LAYER ME3 ;
  RECT 0.000 113.460 1.120 116.700 ;
  LAYER ME2 ;
  RECT 0.000 113.460 1.120 116.700 ;
  LAYER ME1 ;
  RECT 0.000 113.460 1.120 116.700 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 105.620 1.120 108.860 ;
  LAYER ME4 ;
  RECT 0.000 105.620 1.120 108.860 ;
  LAYER ME3 ;
  RECT 0.000 105.620 1.120 108.860 ;
  LAYER ME2 ;
  RECT 0.000 105.620 1.120 108.860 ;
  LAYER ME1 ;
  RECT 0.000 105.620 1.120 108.860 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 97.780 1.120 101.020 ;
  LAYER ME4 ;
  RECT 0.000 97.780 1.120 101.020 ;
  LAYER ME3 ;
  RECT 0.000 97.780 1.120 101.020 ;
  LAYER ME2 ;
  RECT 0.000 97.780 1.120 101.020 ;
  LAYER ME1 ;
  RECT 0.000 97.780 1.120 101.020 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 89.940 1.120 93.180 ;
  LAYER ME4 ;
  RECT 0.000 89.940 1.120 93.180 ;
  LAYER ME3 ;
  RECT 0.000 89.940 1.120 93.180 ;
  LAYER ME2 ;
  RECT 0.000 89.940 1.120 93.180 ;
  LAYER ME1 ;
  RECT 0.000 89.940 1.120 93.180 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 50.740 1.120 53.980 ;
  LAYER ME4 ;
  RECT 0.000 50.740 1.120 53.980 ;
  LAYER ME3 ;
  RECT 0.000 50.740 1.120 53.980 ;
  LAYER ME2 ;
  RECT 0.000 50.740 1.120 53.980 ;
  LAYER ME1 ;
  RECT 0.000 50.740 1.120 53.980 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 42.900 1.120 46.140 ;
  LAYER ME4 ;
  RECT 0.000 42.900 1.120 46.140 ;
  LAYER ME3 ;
  RECT 0.000 42.900 1.120 46.140 ;
  LAYER ME2 ;
  RECT 0.000 42.900 1.120 46.140 ;
  LAYER ME1 ;
  RECT 0.000 42.900 1.120 46.140 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 35.060 1.120 38.300 ;
  LAYER ME4 ;
  RECT 0.000 35.060 1.120 38.300 ;
  LAYER ME3 ;
  RECT 0.000 35.060 1.120 38.300 ;
  LAYER ME2 ;
  RECT 0.000 35.060 1.120 38.300 ;
  LAYER ME1 ;
  RECT 0.000 35.060 1.120 38.300 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 27.220 1.120 30.460 ;
  LAYER ME4 ;
  RECT 0.000 27.220 1.120 30.460 ;
  LAYER ME3 ;
  RECT 0.000 27.220 1.120 30.460 ;
  LAYER ME2 ;
  RECT 0.000 27.220 1.120 30.460 ;
  LAYER ME1 ;
  RECT 0.000 27.220 1.120 30.460 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 19.380 1.120 22.620 ;
  LAYER ME4 ;
  RECT 0.000 19.380 1.120 22.620 ;
  LAYER ME3 ;
  RECT 0.000 19.380 1.120 22.620 ;
  LAYER ME2 ;
  RECT 0.000 19.380 1.120 22.620 ;
  LAYER ME1 ;
  RECT 0.000 19.380 1.120 22.620 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 11.540 1.120 14.780 ;
  LAYER ME4 ;
  RECT 0.000 11.540 1.120 14.780 ;
  LAYER ME3 ;
  RECT 0.000 11.540 1.120 14.780 ;
  LAYER ME2 ;
  RECT 0.000 11.540 1.120 14.780 ;
  LAYER ME1 ;
  RECT 0.000 11.540 1.120 14.780 ;
 END
 PORT
  LAYER ME5 ;
  RECT 911.800 251.440 915.340 252.560 ;
  LAYER ME4 ;
  RECT 911.800 251.440 915.340 252.560 ;
  LAYER ME3 ;
  RECT 911.800 251.440 915.340 252.560 ;
  LAYER ME2 ;
  RECT 911.800 251.440 915.340 252.560 ;
  LAYER ME1 ;
  RECT 911.800 251.440 915.340 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 898.160 251.440 901.700 252.560 ;
  LAYER ME4 ;
  RECT 898.160 251.440 901.700 252.560 ;
  LAYER ME3 ;
  RECT 898.160 251.440 901.700 252.560 ;
  LAYER ME2 ;
  RECT 898.160 251.440 901.700 252.560 ;
  LAYER ME1 ;
  RECT 898.160 251.440 901.700 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 885.140 251.440 888.680 252.560 ;
  LAYER ME4 ;
  RECT 885.140 251.440 888.680 252.560 ;
  LAYER ME3 ;
  RECT 885.140 251.440 888.680 252.560 ;
  LAYER ME2 ;
  RECT 885.140 251.440 888.680 252.560 ;
  LAYER ME1 ;
  RECT 885.140 251.440 888.680 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 871.500 251.440 875.040 252.560 ;
  LAYER ME4 ;
  RECT 871.500 251.440 875.040 252.560 ;
  LAYER ME3 ;
  RECT 871.500 251.440 875.040 252.560 ;
  LAYER ME2 ;
  RECT 871.500 251.440 875.040 252.560 ;
  LAYER ME1 ;
  RECT 871.500 251.440 875.040 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 857.860 251.440 861.400 252.560 ;
  LAYER ME4 ;
  RECT 857.860 251.440 861.400 252.560 ;
  LAYER ME3 ;
  RECT 857.860 251.440 861.400 252.560 ;
  LAYER ME2 ;
  RECT 857.860 251.440 861.400 252.560 ;
  LAYER ME1 ;
  RECT 857.860 251.440 861.400 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 844.840 251.440 848.380 252.560 ;
  LAYER ME4 ;
  RECT 844.840 251.440 848.380 252.560 ;
  LAYER ME3 ;
  RECT 844.840 251.440 848.380 252.560 ;
  LAYER ME2 ;
  RECT 844.840 251.440 848.380 252.560 ;
  LAYER ME1 ;
  RECT 844.840 251.440 848.380 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 777.260 251.440 780.800 252.560 ;
  LAYER ME4 ;
  RECT 777.260 251.440 780.800 252.560 ;
  LAYER ME3 ;
  RECT 777.260 251.440 780.800 252.560 ;
  LAYER ME2 ;
  RECT 777.260 251.440 780.800 252.560 ;
  LAYER ME1 ;
  RECT 777.260 251.440 780.800 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 763.620 251.440 767.160 252.560 ;
  LAYER ME4 ;
  RECT 763.620 251.440 767.160 252.560 ;
  LAYER ME3 ;
  RECT 763.620 251.440 767.160 252.560 ;
  LAYER ME2 ;
  RECT 763.620 251.440 767.160 252.560 ;
  LAYER ME1 ;
  RECT 763.620 251.440 767.160 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 750.600 251.440 754.140 252.560 ;
  LAYER ME4 ;
  RECT 750.600 251.440 754.140 252.560 ;
  LAYER ME3 ;
  RECT 750.600 251.440 754.140 252.560 ;
  LAYER ME2 ;
  RECT 750.600 251.440 754.140 252.560 ;
  LAYER ME1 ;
  RECT 750.600 251.440 754.140 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 736.960 251.440 740.500 252.560 ;
  LAYER ME4 ;
  RECT 736.960 251.440 740.500 252.560 ;
  LAYER ME3 ;
  RECT 736.960 251.440 740.500 252.560 ;
  LAYER ME2 ;
  RECT 736.960 251.440 740.500 252.560 ;
  LAYER ME1 ;
  RECT 736.960 251.440 740.500 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 723.320 251.440 726.860 252.560 ;
  LAYER ME4 ;
  RECT 723.320 251.440 726.860 252.560 ;
  LAYER ME3 ;
  RECT 723.320 251.440 726.860 252.560 ;
  LAYER ME2 ;
  RECT 723.320 251.440 726.860 252.560 ;
  LAYER ME1 ;
  RECT 723.320 251.440 726.860 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 710.300 251.440 713.840 252.560 ;
  LAYER ME4 ;
  RECT 710.300 251.440 713.840 252.560 ;
  LAYER ME3 ;
  RECT 710.300 251.440 713.840 252.560 ;
  LAYER ME2 ;
  RECT 710.300 251.440 713.840 252.560 ;
  LAYER ME1 ;
  RECT 710.300 251.440 713.840 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 642.720 251.440 646.260 252.560 ;
  LAYER ME4 ;
  RECT 642.720 251.440 646.260 252.560 ;
  LAYER ME3 ;
  RECT 642.720 251.440 646.260 252.560 ;
  LAYER ME2 ;
  RECT 642.720 251.440 646.260 252.560 ;
  LAYER ME1 ;
  RECT 642.720 251.440 646.260 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 629.700 251.440 633.240 252.560 ;
  LAYER ME4 ;
  RECT 629.700 251.440 633.240 252.560 ;
  LAYER ME3 ;
  RECT 629.700 251.440 633.240 252.560 ;
  LAYER ME2 ;
  RECT 629.700 251.440 633.240 252.560 ;
  LAYER ME1 ;
  RECT 629.700 251.440 633.240 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 616.060 251.440 619.600 252.560 ;
  LAYER ME4 ;
  RECT 616.060 251.440 619.600 252.560 ;
  LAYER ME3 ;
  RECT 616.060 251.440 619.600 252.560 ;
  LAYER ME2 ;
  RECT 616.060 251.440 619.600 252.560 ;
  LAYER ME1 ;
  RECT 616.060 251.440 619.600 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 602.420 251.440 605.960 252.560 ;
  LAYER ME4 ;
  RECT 602.420 251.440 605.960 252.560 ;
  LAYER ME3 ;
  RECT 602.420 251.440 605.960 252.560 ;
  LAYER ME2 ;
  RECT 602.420 251.440 605.960 252.560 ;
  LAYER ME1 ;
  RECT 602.420 251.440 605.960 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 589.400 251.440 592.940 252.560 ;
  LAYER ME4 ;
  RECT 589.400 251.440 592.940 252.560 ;
  LAYER ME3 ;
  RECT 589.400 251.440 592.940 252.560 ;
  LAYER ME2 ;
  RECT 589.400 251.440 592.940 252.560 ;
  LAYER ME1 ;
  RECT 589.400 251.440 592.940 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 575.760 251.440 579.300 252.560 ;
  LAYER ME4 ;
  RECT 575.760 251.440 579.300 252.560 ;
  LAYER ME3 ;
  RECT 575.760 251.440 579.300 252.560 ;
  LAYER ME2 ;
  RECT 575.760 251.440 579.300 252.560 ;
  LAYER ME1 ;
  RECT 575.760 251.440 579.300 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 513.760 251.440 517.300 252.560 ;
  LAYER ME4 ;
  RECT 513.760 251.440 517.300 252.560 ;
  LAYER ME3 ;
  RECT 513.760 251.440 517.300 252.560 ;
  LAYER ME2 ;
  RECT 513.760 251.440 517.300 252.560 ;
  LAYER ME1 ;
  RECT 513.760 251.440 517.300 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 468.500 251.440 472.040 252.560 ;
  LAYER ME4 ;
  RECT 468.500 251.440 472.040 252.560 ;
  LAYER ME3 ;
  RECT 468.500 251.440 472.040 252.560 ;
  LAYER ME2 ;
  RECT 468.500 251.440 472.040 252.560 ;
  LAYER ME1 ;
  RECT 468.500 251.440 472.040 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 459.820 251.440 463.360 252.560 ;
  LAYER ME4 ;
  RECT 459.820 251.440 463.360 252.560 ;
  LAYER ME3 ;
  RECT 459.820 251.440 463.360 252.560 ;
  LAYER ME2 ;
  RECT 459.820 251.440 463.360 252.560 ;
  LAYER ME1 ;
  RECT 459.820 251.440 463.360 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 439.980 251.440 443.520 252.560 ;
  LAYER ME4 ;
  RECT 439.980 251.440 443.520 252.560 ;
  LAYER ME3 ;
  RECT 439.980 251.440 443.520 252.560 ;
  LAYER ME2 ;
  RECT 439.980 251.440 443.520 252.560 ;
  LAYER ME1 ;
  RECT 439.980 251.440 443.520 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 431.300 251.440 434.840 252.560 ;
  LAYER ME4 ;
  RECT 431.300 251.440 434.840 252.560 ;
  LAYER ME3 ;
  RECT 431.300 251.440 434.840 252.560 ;
  LAYER ME2 ;
  RECT 431.300 251.440 434.840 252.560 ;
  LAYER ME1 ;
  RECT 431.300 251.440 434.840 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 418.280 251.440 421.820 252.560 ;
  LAYER ME4 ;
  RECT 418.280 251.440 421.820 252.560 ;
  LAYER ME3 ;
  RECT 418.280 251.440 421.820 252.560 ;
  LAYER ME2 ;
  RECT 418.280 251.440 421.820 252.560 ;
  LAYER ME1 ;
  RECT 418.280 251.440 421.820 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 350.700 251.440 354.240 252.560 ;
  LAYER ME4 ;
  RECT 350.700 251.440 354.240 252.560 ;
  LAYER ME3 ;
  RECT 350.700 251.440 354.240 252.560 ;
  LAYER ME2 ;
  RECT 350.700 251.440 354.240 252.560 ;
  LAYER ME1 ;
  RECT 350.700 251.440 354.240 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 337.680 251.440 341.220 252.560 ;
  LAYER ME4 ;
  RECT 337.680 251.440 341.220 252.560 ;
  LAYER ME3 ;
  RECT 337.680 251.440 341.220 252.560 ;
  LAYER ME2 ;
  RECT 337.680 251.440 341.220 252.560 ;
  LAYER ME1 ;
  RECT 337.680 251.440 341.220 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 324.040 251.440 327.580 252.560 ;
  LAYER ME4 ;
  RECT 324.040 251.440 327.580 252.560 ;
  LAYER ME3 ;
  RECT 324.040 251.440 327.580 252.560 ;
  LAYER ME2 ;
  RECT 324.040 251.440 327.580 252.560 ;
  LAYER ME1 ;
  RECT 324.040 251.440 327.580 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 310.400 251.440 313.940 252.560 ;
  LAYER ME4 ;
  RECT 310.400 251.440 313.940 252.560 ;
  LAYER ME3 ;
  RECT 310.400 251.440 313.940 252.560 ;
  LAYER ME2 ;
  RECT 310.400 251.440 313.940 252.560 ;
  LAYER ME1 ;
  RECT 310.400 251.440 313.940 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 297.380 251.440 300.920 252.560 ;
  LAYER ME4 ;
  RECT 297.380 251.440 300.920 252.560 ;
  LAYER ME3 ;
  RECT 297.380 251.440 300.920 252.560 ;
  LAYER ME2 ;
  RECT 297.380 251.440 300.920 252.560 ;
  LAYER ME1 ;
  RECT 297.380 251.440 300.920 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 283.740 251.440 287.280 252.560 ;
  LAYER ME4 ;
  RECT 283.740 251.440 287.280 252.560 ;
  LAYER ME3 ;
  RECT 283.740 251.440 287.280 252.560 ;
  LAYER ME2 ;
  RECT 283.740 251.440 287.280 252.560 ;
  LAYER ME1 ;
  RECT 283.740 251.440 287.280 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 216.780 251.440 220.320 252.560 ;
  LAYER ME4 ;
  RECT 216.780 251.440 220.320 252.560 ;
  LAYER ME3 ;
  RECT 216.780 251.440 220.320 252.560 ;
  LAYER ME2 ;
  RECT 216.780 251.440 220.320 252.560 ;
  LAYER ME1 ;
  RECT 216.780 251.440 220.320 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 203.140 251.440 206.680 252.560 ;
  LAYER ME4 ;
  RECT 203.140 251.440 206.680 252.560 ;
  LAYER ME3 ;
  RECT 203.140 251.440 206.680 252.560 ;
  LAYER ME2 ;
  RECT 203.140 251.440 206.680 252.560 ;
  LAYER ME1 ;
  RECT 203.140 251.440 206.680 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 189.500 251.440 193.040 252.560 ;
  LAYER ME4 ;
  RECT 189.500 251.440 193.040 252.560 ;
  LAYER ME3 ;
  RECT 189.500 251.440 193.040 252.560 ;
  LAYER ME2 ;
  RECT 189.500 251.440 193.040 252.560 ;
  LAYER ME1 ;
  RECT 189.500 251.440 193.040 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 176.480 251.440 180.020 252.560 ;
  LAYER ME4 ;
  RECT 176.480 251.440 180.020 252.560 ;
  LAYER ME3 ;
  RECT 176.480 251.440 180.020 252.560 ;
  LAYER ME2 ;
  RECT 176.480 251.440 180.020 252.560 ;
  LAYER ME1 ;
  RECT 176.480 251.440 180.020 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 162.840 251.440 166.380 252.560 ;
  LAYER ME4 ;
  RECT 162.840 251.440 166.380 252.560 ;
  LAYER ME3 ;
  RECT 162.840 251.440 166.380 252.560 ;
  LAYER ME2 ;
  RECT 162.840 251.440 166.380 252.560 ;
  LAYER ME1 ;
  RECT 162.840 251.440 166.380 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 149.200 251.440 152.740 252.560 ;
  LAYER ME4 ;
  RECT 149.200 251.440 152.740 252.560 ;
  LAYER ME3 ;
  RECT 149.200 251.440 152.740 252.560 ;
  LAYER ME2 ;
  RECT 149.200 251.440 152.740 252.560 ;
  LAYER ME1 ;
  RECT 149.200 251.440 152.740 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 82.240 251.440 85.780 252.560 ;
  LAYER ME4 ;
  RECT 82.240 251.440 85.780 252.560 ;
  LAYER ME3 ;
  RECT 82.240 251.440 85.780 252.560 ;
  LAYER ME2 ;
  RECT 82.240 251.440 85.780 252.560 ;
  LAYER ME1 ;
  RECT 82.240 251.440 85.780 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 68.600 251.440 72.140 252.560 ;
  LAYER ME4 ;
  RECT 68.600 251.440 72.140 252.560 ;
  LAYER ME3 ;
  RECT 68.600 251.440 72.140 252.560 ;
  LAYER ME2 ;
  RECT 68.600 251.440 72.140 252.560 ;
  LAYER ME1 ;
  RECT 68.600 251.440 72.140 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 54.960 251.440 58.500 252.560 ;
  LAYER ME4 ;
  RECT 54.960 251.440 58.500 252.560 ;
  LAYER ME3 ;
  RECT 54.960 251.440 58.500 252.560 ;
  LAYER ME2 ;
  RECT 54.960 251.440 58.500 252.560 ;
  LAYER ME1 ;
  RECT 54.960 251.440 58.500 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 41.940 251.440 45.480 252.560 ;
  LAYER ME4 ;
  RECT 41.940 251.440 45.480 252.560 ;
  LAYER ME3 ;
  RECT 41.940 251.440 45.480 252.560 ;
  LAYER ME2 ;
  RECT 41.940 251.440 45.480 252.560 ;
  LAYER ME1 ;
  RECT 41.940 251.440 45.480 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 28.300 251.440 31.840 252.560 ;
  LAYER ME4 ;
  RECT 28.300 251.440 31.840 252.560 ;
  LAYER ME3 ;
  RECT 28.300 251.440 31.840 252.560 ;
  LAYER ME2 ;
  RECT 28.300 251.440 31.840 252.560 ;
  LAYER ME1 ;
  RECT 28.300 251.440 31.840 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 14.660 251.440 18.200 252.560 ;
  LAYER ME4 ;
  RECT 14.660 251.440 18.200 252.560 ;
  LAYER ME3 ;
  RECT 14.660 251.440 18.200 252.560 ;
  LAYER ME2 ;
  RECT 14.660 251.440 18.200 252.560 ;
  LAYER ME1 ;
  RECT 14.660 251.440 18.200 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 911.800 0.000 915.340 1.120 ;
  LAYER ME4 ;
  RECT 911.800 0.000 915.340 1.120 ;
  LAYER ME3 ;
  RECT 911.800 0.000 915.340 1.120 ;
  LAYER ME2 ;
  RECT 911.800 0.000 915.340 1.120 ;
  LAYER ME1 ;
  RECT 911.800 0.000 915.340 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 898.160 0.000 901.700 1.120 ;
  LAYER ME4 ;
  RECT 898.160 0.000 901.700 1.120 ;
  LAYER ME3 ;
  RECT 898.160 0.000 901.700 1.120 ;
  LAYER ME2 ;
  RECT 898.160 0.000 901.700 1.120 ;
  LAYER ME1 ;
  RECT 898.160 0.000 901.700 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 885.140 0.000 888.680 1.120 ;
  LAYER ME4 ;
  RECT 885.140 0.000 888.680 1.120 ;
  LAYER ME3 ;
  RECT 885.140 0.000 888.680 1.120 ;
  LAYER ME2 ;
  RECT 885.140 0.000 888.680 1.120 ;
  LAYER ME1 ;
  RECT 885.140 0.000 888.680 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 871.500 0.000 875.040 1.120 ;
  LAYER ME4 ;
  RECT 871.500 0.000 875.040 1.120 ;
  LAYER ME3 ;
  RECT 871.500 0.000 875.040 1.120 ;
  LAYER ME2 ;
  RECT 871.500 0.000 875.040 1.120 ;
  LAYER ME1 ;
  RECT 871.500 0.000 875.040 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 857.860 0.000 861.400 1.120 ;
  LAYER ME4 ;
  RECT 857.860 0.000 861.400 1.120 ;
  LAYER ME3 ;
  RECT 857.860 0.000 861.400 1.120 ;
  LAYER ME2 ;
  RECT 857.860 0.000 861.400 1.120 ;
  LAYER ME1 ;
  RECT 857.860 0.000 861.400 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 844.840 0.000 848.380 1.120 ;
  LAYER ME4 ;
  RECT 844.840 0.000 848.380 1.120 ;
  LAYER ME3 ;
  RECT 844.840 0.000 848.380 1.120 ;
  LAYER ME2 ;
  RECT 844.840 0.000 848.380 1.120 ;
  LAYER ME1 ;
  RECT 844.840 0.000 848.380 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 777.260 0.000 780.800 1.120 ;
  LAYER ME4 ;
  RECT 777.260 0.000 780.800 1.120 ;
  LAYER ME3 ;
  RECT 777.260 0.000 780.800 1.120 ;
  LAYER ME2 ;
  RECT 777.260 0.000 780.800 1.120 ;
  LAYER ME1 ;
  RECT 777.260 0.000 780.800 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 763.620 0.000 767.160 1.120 ;
  LAYER ME4 ;
  RECT 763.620 0.000 767.160 1.120 ;
  LAYER ME3 ;
  RECT 763.620 0.000 767.160 1.120 ;
  LAYER ME2 ;
  RECT 763.620 0.000 767.160 1.120 ;
  LAYER ME1 ;
  RECT 763.620 0.000 767.160 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 750.600 0.000 754.140 1.120 ;
  LAYER ME4 ;
  RECT 750.600 0.000 754.140 1.120 ;
  LAYER ME3 ;
  RECT 750.600 0.000 754.140 1.120 ;
  LAYER ME2 ;
  RECT 750.600 0.000 754.140 1.120 ;
  LAYER ME1 ;
  RECT 750.600 0.000 754.140 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 736.960 0.000 740.500 1.120 ;
  LAYER ME4 ;
  RECT 736.960 0.000 740.500 1.120 ;
  LAYER ME3 ;
  RECT 736.960 0.000 740.500 1.120 ;
  LAYER ME2 ;
  RECT 736.960 0.000 740.500 1.120 ;
  LAYER ME1 ;
  RECT 736.960 0.000 740.500 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 723.320 0.000 726.860 1.120 ;
  LAYER ME4 ;
  RECT 723.320 0.000 726.860 1.120 ;
  LAYER ME3 ;
  RECT 723.320 0.000 726.860 1.120 ;
  LAYER ME2 ;
  RECT 723.320 0.000 726.860 1.120 ;
  LAYER ME1 ;
  RECT 723.320 0.000 726.860 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 710.300 0.000 713.840 1.120 ;
  LAYER ME4 ;
  RECT 710.300 0.000 713.840 1.120 ;
  LAYER ME3 ;
  RECT 710.300 0.000 713.840 1.120 ;
  LAYER ME2 ;
  RECT 710.300 0.000 713.840 1.120 ;
  LAYER ME1 ;
  RECT 710.300 0.000 713.840 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 642.720 0.000 646.260 1.120 ;
  LAYER ME4 ;
  RECT 642.720 0.000 646.260 1.120 ;
  LAYER ME3 ;
  RECT 642.720 0.000 646.260 1.120 ;
  LAYER ME2 ;
  RECT 642.720 0.000 646.260 1.120 ;
  LAYER ME1 ;
  RECT 642.720 0.000 646.260 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 629.700 0.000 633.240 1.120 ;
  LAYER ME4 ;
  RECT 629.700 0.000 633.240 1.120 ;
  LAYER ME3 ;
  RECT 629.700 0.000 633.240 1.120 ;
  LAYER ME2 ;
  RECT 629.700 0.000 633.240 1.120 ;
  LAYER ME1 ;
  RECT 629.700 0.000 633.240 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 616.060 0.000 619.600 1.120 ;
  LAYER ME4 ;
  RECT 616.060 0.000 619.600 1.120 ;
  LAYER ME3 ;
  RECT 616.060 0.000 619.600 1.120 ;
  LAYER ME2 ;
  RECT 616.060 0.000 619.600 1.120 ;
  LAYER ME1 ;
  RECT 616.060 0.000 619.600 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 602.420 0.000 605.960 1.120 ;
  LAYER ME4 ;
  RECT 602.420 0.000 605.960 1.120 ;
  LAYER ME3 ;
  RECT 602.420 0.000 605.960 1.120 ;
  LAYER ME2 ;
  RECT 602.420 0.000 605.960 1.120 ;
  LAYER ME1 ;
  RECT 602.420 0.000 605.960 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 589.400 0.000 592.940 1.120 ;
  LAYER ME4 ;
  RECT 589.400 0.000 592.940 1.120 ;
  LAYER ME3 ;
  RECT 589.400 0.000 592.940 1.120 ;
  LAYER ME2 ;
  RECT 589.400 0.000 592.940 1.120 ;
  LAYER ME1 ;
  RECT 589.400 0.000 592.940 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 575.760 0.000 579.300 1.120 ;
  LAYER ME4 ;
  RECT 575.760 0.000 579.300 1.120 ;
  LAYER ME3 ;
  RECT 575.760 0.000 579.300 1.120 ;
  LAYER ME2 ;
  RECT 575.760 0.000 579.300 1.120 ;
  LAYER ME1 ;
  RECT 575.760 0.000 579.300 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 513.760 0.000 517.300 1.120 ;
  LAYER ME4 ;
  RECT 513.760 0.000 517.300 1.120 ;
  LAYER ME3 ;
  RECT 513.760 0.000 517.300 1.120 ;
  LAYER ME2 ;
  RECT 513.760 0.000 517.300 1.120 ;
  LAYER ME1 ;
  RECT 513.760 0.000 517.300 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 468.500 0.000 472.040 1.120 ;
  LAYER ME4 ;
  RECT 468.500 0.000 472.040 1.120 ;
  LAYER ME3 ;
  RECT 468.500 0.000 472.040 1.120 ;
  LAYER ME2 ;
  RECT 468.500 0.000 472.040 1.120 ;
  LAYER ME1 ;
  RECT 468.500 0.000 472.040 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 459.820 0.000 463.360 1.120 ;
  LAYER ME4 ;
  RECT 459.820 0.000 463.360 1.120 ;
  LAYER ME3 ;
  RECT 459.820 0.000 463.360 1.120 ;
  LAYER ME2 ;
  RECT 459.820 0.000 463.360 1.120 ;
  LAYER ME1 ;
  RECT 459.820 0.000 463.360 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 439.980 0.000 443.520 1.120 ;
  LAYER ME4 ;
  RECT 439.980 0.000 443.520 1.120 ;
  LAYER ME3 ;
  RECT 439.980 0.000 443.520 1.120 ;
  LAYER ME2 ;
  RECT 439.980 0.000 443.520 1.120 ;
  LAYER ME1 ;
  RECT 439.980 0.000 443.520 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 431.300 0.000 434.840 1.120 ;
  LAYER ME4 ;
  RECT 431.300 0.000 434.840 1.120 ;
  LAYER ME3 ;
  RECT 431.300 0.000 434.840 1.120 ;
  LAYER ME2 ;
  RECT 431.300 0.000 434.840 1.120 ;
  LAYER ME1 ;
  RECT 431.300 0.000 434.840 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 418.280 0.000 421.820 1.120 ;
  LAYER ME4 ;
  RECT 418.280 0.000 421.820 1.120 ;
  LAYER ME3 ;
  RECT 418.280 0.000 421.820 1.120 ;
  LAYER ME2 ;
  RECT 418.280 0.000 421.820 1.120 ;
  LAYER ME1 ;
  RECT 418.280 0.000 421.820 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 350.700 0.000 354.240 1.120 ;
  LAYER ME4 ;
  RECT 350.700 0.000 354.240 1.120 ;
  LAYER ME3 ;
  RECT 350.700 0.000 354.240 1.120 ;
  LAYER ME2 ;
  RECT 350.700 0.000 354.240 1.120 ;
  LAYER ME1 ;
  RECT 350.700 0.000 354.240 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 337.680 0.000 341.220 1.120 ;
  LAYER ME4 ;
  RECT 337.680 0.000 341.220 1.120 ;
  LAYER ME3 ;
  RECT 337.680 0.000 341.220 1.120 ;
  LAYER ME2 ;
  RECT 337.680 0.000 341.220 1.120 ;
  LAYER ME1 ;
  RECT 337.680 0.000 341.220 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 324.040 0.000 327.580 1.120 ;
  LAYER ME4 ;
  RECT 324.040 0.000 327.580 1.120 ;
  LAYER ME3 ;
  RECT 324.040 0.000 327.580 1.120 ;
  LAYER ME2 ;
  RECT 324.040 0.000 327.580 1.120 ;
  LAYER ME1 ;
  RECT 324.040 0.000 327.580 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 310.400 0.000 313.940 1.120 ;
  LAYER ME4 ;
  RECT 310.400 0.000 313.940 1.120 ;
  LAYER ME3 ;
  RECT 310.400 0.000 313.940 1.120 ;
  LAYER ME2 ;
  RECT 310.400 0.000 313.940 1.120 ;
  LAYER ME1 ;
  RECT 310.400 0.000 313.940 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 297.380 0.000 300.920 1.120 ;
  LAYER ME4 ;
  RECT 297.380 0.000 300.920 1.120 ;
  LAYER ME3 ;
  RECT 297.380 0.000 300.920 1.120 ;
  LAYER ME2 ;
  RECT 297.380 0.000 300.920 1.120 ;
  LAYER ME1 ;
  RECT 297.380 0.000 300.920 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 283.740 0.000 287.280 1.120 ;
  LAYER ME4 ;
  RECT 283.740 0.000 287.280 1.120 ;
  LAYER ME3 ;
  RECT 283.740 0.000 287.280 1.120 ;
  LAYER ME2 ;
  RECT 283.740 0.000 287.280 1.120 ;
  LAYER ME1 ;
  RECT 283.740 0.000 287.280 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 216.780 0.000 220.320 1.120 ;
  LAYER ME4 ;
  RECT 216.780 0.000 220.320 1.120 ;
  LAYER ME3 ;
  RECT 216.780 0.000 220.320 1.120 ;
  LAYER ME2 ;
  RECT 216.780 0.000 220.320 1.120 ;
  LAYER ME1 ;
  RECT 216.780 0.000 220.320 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 203.140 0.000 206.680 1.120 ;
  LAYER ME4 ;
  RECT 203.140 0.000 206.680 1.120 ;
  LAYER ME3 ;
  RECT 203.140 0.000 206.680 1.120 ;
  LAYER ME2 ;
  RECT 203.140 0.000 206.680 1.120 ;
  LAYER ME1 ;
  RECT 203.140 0.000 206.680 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 189.500 0.000 193.040 1.120 ;
  LAYER ME4 ;
  RECT 189.500 0.000 193.040 1.120 ;
  LAYER ME3 ;
  RECT 189.500 0.000 193.040 1.120 ;
  LAYER ME2 ;
  RECT 189.500 0.000 193.040 1.120 ;
  LAYER ME1 ;
  RECT 189.500 0.000 193.040 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 176.480 0.000 180.020 1.120 ;
  LAYER ME4 ;
  RECT 176.480 0.000 180.020 1.120 ;
  LAYER ME3 ;
  RECT 176.480 0.000 180.020 1.120 ;
  LAYER ME2 ;
  RECT 176.480 0.000 180.020 1.120 ;
  LAYER ME1 ;
  RECT 176.480 0.000 180.020 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 162.840 0.000 166.380 1.120 ;
  LAYER ME4 ;
  RECT 162.840 0.000 166.380 1.120 ;
  LAYER ME3 ;
  RECT 162.840 0.000 166.380 1.120 ;
  LAYER ME2 ;
  RECT 162.840 0.000 166.380 1.120 ;
  LAYER ME1 ;
  RECT 162.840 0.000 166.380 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 149.200 0.000 152.740 1.120 ;
  LAYER ME4 ;
  RECT 149.200 0.000 152.740 1.120 ;
  LAYER ME3 ;
  RECT 149.200 0.000 152.740 1.120 ;
  LAYER ME2 ;
  RECT 149.200 0.000 152.740 1.120 ;
  LAYER ME1 ;
  RECT 149.200 0.000 152.740 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 82.240 0.000 85.780 1.120 ;
  LAYER ME4 ;
  RECT 82.240 0.000 85.780 1.120 ;
  LAYER ME3 ;
  RECT 82.240 0.000 85.780 1.120 ;
  LAYER ME2 ;
  RECT 82.240 0.000 85.780 1.120 ;
  LAYER ME1 ;
  RECT 82.240 0.000 85.780 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 68.600 0.000 72.140 1.120 ;
  LAYER ME4 ;
  RECT 68.600 0.000 72.140 1.120 ;
  LAYER ME3 ;
  RECT 68.600 0.000 72.140 1.120 ;
  LAYER ME2 ;
  RECT 68.600 0.000 72.140 1.120 ;
  LAYER ME1 ;
  RECT 68.600 0.000 72.140 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 54.960 0.000 58.500 1.120 ;
  LAYER ME4 ;
  RECT 54.960 0.000 58.500 1.120 ;
  LAYER ME3 ;
  RECT 54.960 0.000 58.500 1.120 ;
  LAYER ME2 ;
  RECT 54.960 0.000 58.500 1.120 ;
  LAYER ME1 ;
  RECT 54.960 0.000 58.500 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 41.940 0.000 45.480 1.120 ;
  LAYER ME4 ;
  RECT 41.940 0.000 45.480 1.120 ;
  LAYER ME3 ;
  RECT 41.940 0.000 45.480 1.120 ;
  LAYER ME2 ;
  RECT 41.940 0.000 45.480 1.120 ;
  LAYER ME1 ;
  RECT 41.940 0.000 45.480 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 28.300 0.000 31.840 1.120 ;
  LAYER ME4 ;
  RECT 28.300 0.000 31.840 1.120 ;
  LAYER ME3 ;
  RECT 28.300 0.000 31.840 1.120 ;
  LAYER ME2 ;
  RECT 28.300 0.000 31.840 1.120 ;
  LAYER ME1 ;
  RECT 28.300 0.000 31.840 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 14.660 0.000 18.200 1.120 ;
  LAYER ME4 ;
  RECT 14.660 0.000 18.200 1.120 ;
  LAYER ME3 ;
  RECT 14.660 0.000 18.200 1.120 ;
  LAYER ME2 ;
  RECT 14.660 0.000 18.200 1.120 ;
  LAYER ME1 ;
  RECT 14.660 0.000 18.200 1.120 ;
 END
END GND
PIN VCC
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
 PORT
  LAYER ME5 ;
  RECT 971.660 203.620 972.780 206.860 ;
  LAYER ME4 ;
  RECT 971.660 203.620 972.780 206.860 ;
  LAYER ME3 ;
  RECT 971.660 203.620 972.780 206.860 ;
  LAYER ME2 ;
  RECT 971.660 203.620 972.780 206.860 ;
  LAYER ME1 ;
  RECT 971.660 203.620 972.780 206.860 ;
 END
 PORT
  LAYER ME5 ;
  RECT 971.660 195.780 972.780 199.020 ;
  LAYER ME4 ;
  RECT 971.660 195.780 972.780 199.020 ;
  LAYER ME3 ;
  RECT 971.660 195.780 972.780 199.020 ;
  LAYER ME2 ;
  RECT 971.660 195.780 972.780 199.020 ;
  LAYER ME1 ;
  RECT 971.660 195.780 972.780 199.020 ;
 END
 PORT
  LAYER ME5 ;
  RECT 971.660 187.940 972.780 191.180 ;
  LAYER ME4 ;
  RECT 971.660 187.940 972.780 191.180 ;
  LAYER ME3 ;
  RECT 971.660 187.940 972.780 191.180 ;
  LAYER ME2 ;
  RECT 971.660 187.940 972.780 191.180 ;
  LAYER ME1 ;
  RECT 971.660 187.940 972.780 191.180 ;
 END
 PORT
  LAYER ME5 ;
  RECT 971.660 180.100 972.780 183.340 ;
  LAYER ME4 ;
  RECT 971.660 180.100 972.780 183.340 ;
  LAYER ME3 ;
  RECT 971.660 180.100 972.780 183.340 ;
  LAYER ME2 ;
  RECT 971.660 180.100 972.780 183.340 ;
  LAYER ME1 ;
  RECT 971.660 180.100 972.780 183.340 ;
 END
 PORT
  LAYER ME5 ;
  RECT 971.660 172.260 972.780 175.500 ;
  LAYER ME4 ;
  RECT 971.660 172.260 972.780 175.500 ;
  LAYER ME3 ;
  RECT 971.660 172.260 972.780 175.500 ;
  LAYER ME2 ;
  RECT 971.660 172.260 972.780 175.500 ;
  LAYER ME1 ;
  RECT 971.660 172.260 972.780 175.500 ;
 END
 PORT
  LAYER ME5 ;
  RECT 971.660 164.420 972.780 167.660 ;
  LAYER ME4 ;
  RECT 971.660 164.420 972.780 167.660 ;
  LAYER ME3 ;
  RECT 971.660 164.420 972.780 167.660 ;
  LAYER ME2 ;
  RECT 971.660 164.420 972.780 167.660 ;
  LAYER ME1 ;
  RECT 971.660 164.420 972.780 167.660 ;
 END
 PORT
  LAYER ME5 ;
  RECT 971.660 125.220 972.780 128.460 ;
  LAYER ME4 ;
  RECT 971.660 125.220 972.780 128.460 ;
  LAYER ME3 ;
  RECT 971.660 125.220 972.780 128.460 ;
  LAYER ME2 ;
  RECT 971.660 125.220 972.780 128.460 ;
  LAYER ME1 ;
  RECT 971.660 125.220 972.780 128.460 ;
 END
 PORT
  LAYER ME5 ;
  RECT 971.660 117.380 972.780 120.620 ;
  LAYER ME4 ;
  RECT 971.660 117.380 972.780 120.620 ;
  LAYER ME3 ;
  RECT 971.660 117.380 972.780 120.620 ;
  LAYER ME2 ;
  RECT 971.660 117.380 972.780 120.620 ;
  LAYER ME1 ;
  RECT 971.660 117.380 972.780 120.620 ;
 END
 PORT
  LAYER ME5 ;
  RECT 971.660 109.540 972.780 112.780 ;
  LAYER ME4 ;
  RECT 971.660 109.540 972.780 112.780 ;
  LAYER ME3 ;
  RECT 971.660 109.540 972.780 112.780 ;
  LAYER ME2 ;
  RECT 971.660 109.540 972.780 112.780 ;
  LAYER ME1 ;
  RECT 971.660 109.540 972.780 112.780 ;
 END
 PORT
  LAYER ME5 ;
  RECT 971.660 101.700 972.780 104.940 ;
  LAYER ME4 ;
  RECT 971.660 101.700 972.780 104.940 ;
  LAYER ME3 ;
  RECT 971.660 101.700 972.780 104.940 ;
  LAYER ME2 ;
  RECT 971.660 101.700 972.780 104.940 ;
  LAYER ME1 ;
  RECT 971.660 101.700 972.780 104.940 ;
 END
 PORT
  LAYER ME5 ;
  RECT 971.660 93.860 972.780 97.100 ;
  LAYER ME4 ;
  RECT 971.660 93.860 972.780 97.100 ;
  LAYER ME3 ;
  RECT 971.660 93.860 972.780 97.100 ;
  LAYER ME2 ;
  RECT 971.660 93.860 972.780 97.100 ;
  LAYER ME1 ;
  RECT 971.660 93.860 972.780 97.100 ;
 END
 PORT
  LAYER ME5 ;
  RECT 971.660 86.020 972.780 89.260 ;
  LAYER ME4 ;
  RECT 971.660 86.020 972.780 89.260 ;
  LAYER ME3 ;
  RECT 971.660 86.020 972.780 89.260 ;
  LAYER ME2 ;
  RECT 971.660 86.020 972.780 89.260 ;
  LAYER ME1 ;
  RECT 971.660 86.020 972.780 89.260 ;
 END
 PORT
  LAYER ME5 ;
  RECT 971.660 46.820 972.780 50.060 ;
  LAYER ME4 ;
  RECT 971.660 46.820 972.780 50.060 ;
  LAYER ME3 ;
  RECT 971.660 46.820 972.780 50.060 ;
  LAYER ME2 ;
  RECT 971.660 46.820 972.780 50.060 ;
  LAYER ME1 ;
  RECT 971.660 46.820 972.780 50.060 ;
 END
 PORT
  LAYER ME5 ;
  RECT 971.660 38.980 972.780 42.220 ;
  LAYER ME4 ;
  RECT 971.660 38.980 972.780 42.220 ;
  LAYER ME3 ;
  RECT 971.660 38.980 972.780 42.220 ;
  LAYER ME2 ;
  RECT 971.660 38.980 972.780 42.220 ;
  LAYER ME1 ;
  RECT 971.660 38.980 972.780 42.220 ;
 END
 PORT
  LAYER ME5 ;
  RECT 971.660 31.140 972.780 34.380 ;
  LAYER ME4 ;
  RECT 971.660 31.140 972.780 34.380 ;
  LAYER ME3 ;
  RECT 971.660 31.140 972.780 34.380 ;
  LAYER ME2 ;
  RECT 971.660 31.140 972.780 34.380 ;
  LAYER ME1 ;
  RECT 971.660 31.140 972.780 34.380 ;
 END
 PORT
  LAYER ME5 ;
  RECT 971.660 23.300 972.780 26.540 ;
  LAYER ME4 ;
  RECT 971.660 23.300 972.780 26.540 ;
  LAYER ME3 ;
  RECT 971.660 23.300 972.780 26.540 ;
  LAYER ME2 ;
  RECT 971.660 23.300 972.780 26.540 ;
  LAYER ME1 ;
  RECT 971.660 23.300 972.780 26.540 ;
 END
 PORT
  LAYER ME5 ;
  RECT 971.660 15.460 972.780 18.700 ;
  LAYER ME4 ;
  RECT 971.660 15.460 972.780 18.700 ;
  LAYER ME3 ;
  RECT 971.660 15.460 972.780 18.700 ;
  LAYER ME2 ;
  RECT 971.660 15.460 972.780 18.700 ;
  LAYER ME1 ;
  RECT 971.660 15.460 972.780 18.700 ;
 END
 PORT
  LAYER ME5 ;
  RECT 971.660 7.620 972.780 10.860 ;
  LAYER ME4 ;
  RECT 971.660 7.620 972.780 10.860 ;
  LAYER ME3 ;
  RECT 971.660 7.620 972.780 10.860 ;
  LAYER ME2 ;
  RECT 971.660 7.620 972.780 10.860 ;
  LAYER ME1 ;
  RECT 971.660 7.620 972.780 10.860 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 203.620 1.120 206.860 ;
  LAYER ME4 ;
  RECT 0.000 203.620 1.120 206.860 ;
  LAYER ME3 ;
  RECT 0.000 203.620 1.120 206.860 ;
  LAYER ME2 ;
  RECT 0.000 203.620 1.120 206.860 ;
  LAYER ME1 ;
  RECT 0.000 203.620 1.120 206.860 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 195.780 1.120 199.020 ;
  LAYER ME4 ;
  RECT 0.000 195.780 1.120 199.020 ;
  LAYER ME3 ;
  RECT 0.000 195.780 1.120 199.020 ;
  LAYER ME2 ;
  RECT 0.000 195.780 1.120 199.020 ;
  LAYER ME1 ;
  RECT 0.000 195.780 1.120 199.020 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 187.940 1.120 191.180 ;
  LAYER ME4 ;
  RECT 0.000 187.940 1.120 191.180 ;
  LAYER ME3 ;
  RECT 0.000 187.940 1.120 191.180 ;
  LAYER ME2 ;
  RECT 0.000 187.940 1.120 191.180 ;
  LAYER ME1 ;
  RECT 0.000 187.940 1.120 191.180 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 180.100 1.120 183.340 ;
  LAYER ME4 ;
  RECT 0.000 180.100 1.120 183.340 ;
  LAYER ME3 ;
  RECT 0.000 180.100 1.120 183.340 ;
  LAYER ME2 ;
  RECT 0.000 180.100 1.120 183.340 ;
  LAYER ME1 ;
  RECT 0.000 180.100 1.120 183.340 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 172.260 1.120 175.500 ;
  LAYER ME4 ;
  RECT 0.000 172.260 1.120 175.500 ;
  LAYER ME3 ;
  RECT 0.000 172.260 1.120 175.500 ;
  LAYER ME2 ;
  RECT 0.000 172.260 1.120 175.500 ;
  LAYER ME1 ;
  RECT 0.000 172.260 1.120 175.500 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 164.420 1.120 167.660 ;
  LAYER ME4 ;
  RECT 0.000 164.420 1.120 167.660 ;
  LAYER ME3 ;
  RECT 0.000 164.420 1.120 167.660 ;
  LAYER ME2 ;
  RECT 0.000 164.420 1.120 167.660 ;
  LAYER ME1 ;
  RECT 0.000 164.420 1.120 167.660 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 125.220 1.120 128.460 ;
  LAYER ME4 ;
  RECT 0.000 125.220 1.120 128.460 ;
  LAYER ME3 ;
  RECT 0.000 125.220 1.120 128.460 ;
  LAYER ME2 ;
  RECT 0.000 125.220 1.120 128.460 ;
  LAYER ME1 ;
  RECT 0.000 125.220 1.120 128.460 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 117.380 1.120 120.620 ;
  LAYER ME4 ;
  RECT 0.000 117.380 1.120 120.620 ;
  LAYER ME3 ;
  RECT 0.000 117.380 1.120 120.620 ;
  LAYER ME2 ;
  RECT 0.000 117.380 1.120 120.620 ;
  LAYER ME1 ;
  RECT 0.000 117.380 1.120 120.620 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 109.540 1.120 112.780 ;
  LAYER ME4 ;
  RECT 0.000 109.540 1.120 112.780 ;
  LAYER ME3 ;
  RECT 0.000 109.540 1.120 112.780 ;
  LAYER ME2 ;
  RECT 0.000 109.540 1.120 112.780 ;
  LAYER ME1 ;
  RECT 0.000 109.540 1.120 112.780 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 101.700 1.120 104.940 ;
  LAYER ME4 ;
  RECT 0.000 101.700 1.120 104.940 ;
  LAYER ME3 ;
  RECT 0.000 101.700 1.120 104.940 ;
  LAYER ME2 ;
  RECT 0.000 101.700 1.120 104.940 ;
  LAYER ME1 ;
  RECT 0.000 101.700 1.120 104.940 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 93.860 1.120 97.100 ;
  LAYER ME4 ;
  RECT 0.000 93.860 1.120 97.100 ;
  LAYER ME3 ;
  RECT 0.000 93.860 1.120 97.100 ;
  LAYER ME2 ;
  RECT 0.000 93.860 1.120 97.100 ;
  LAYER ME1 ;
  RECT 0.000 93.860 1.120 97.100 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 86.020 1.120 89.260 ;
  LAYER ME4 ;
  RECT 0.000 86.020 1.120 89.260 ;
  LAYER ME3 ;
  RECT 0.000 86.020 1.120 89.260 ;
  LAYER ME2 ;
  RECT 0.000 86.020 1.120 89.260 ;
  LAYER ME1 ;
  RECT 0.000 86.020 1.120 89.260 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 46.820 1.120 50.060 ;
  LAYER ME4 ;
  RECT 0.000 46.820 1.120 50.060 ;
  LAYER ME3 ;
  RECT 0.000 46.820 1.120 50.060 ;
  LAYER ME2 ;
  RECT 0.000 46.820 1.120 50.060 ;
  LAYER ME1 ;
  RECT 0.000 46.820 1.120 50.060 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 38.980 1.120 42.220 ;
  LAYER ME4 ;
  RECT 0.000 38.980 1.120 42.220 ;
  LAYER ME3 ;
  RECT 0.000 38.980 1.120 42.220 ;
  LAYER ME2 ;
  RECT 0.000 38.980 1.120 42.220 ;
  LAYER ME1 ;
  RECT 0.000 38.980 1.120 42.220 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 31.140 1.120 34.380 ;
  LAYER ME4 ;
  RECT 0.000 31.140 1.120 34.380 ;
  LAYER ME3 ;
  RECT 0.000 31.140 1.120 34.380 ;
  LAYER ME2 ;
  RECT 0.000 31.140 1.120 34.380 ;
  LAYER ME1 ;
  RECT 0.000 31.140 1.120 34.380 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 23.300 1.120 26.540 ;
  LAYER ME4 ;
  RECT 0.000 23.300 1.120 26.540 ;
  LAYER ME3 ;
  RECT 0.000 23.300 1.120 26.540 ;
  LAYER ME2 ;
  RECT 0.000 23.300 1.120 26.540 ;
  LAYER ME1 ;
  RECT 0.000 23.300 1.120 26.540 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 15.460 1.120 18.700 ;
  LAYER ME4 ;
  RECT 0.000 15.460 1.120 18.700 ;
  LAYER ME3 ;
  RECT 0.000 15.460 1.120 18.700 ;
  LAYER ME2 ;
  RECT 0.000 15.460 1.120 18.700 ;
  LAYER ME1 ;
  RECT 0.000 15.460 1.120 18.700 ;
 END
 PORT
  LAYER ME5 ;
  RECT 0.000 7.620 1.120 10.860 ;
  LAYER ME4 ;
  RECT 0.000 7.620 1.120 10.860 ;
  LAYER ME3 ;
  RECT 0.000 7.620 1.120 10.860 ;
  LAYER ME2 ;
  RECT 0.000 7.620 1.120 10.860 ;
  LAYER ME1 ;
  RECT 0.000 7.620 1.120 10.860 ;
 END
 PORT
  LAYER ME5 ;
  RECT 902.500 251.440 906.040 252.560 ;
  LAYER ME4 ;
  RECT 902.500 251.440 906.040 252.560 ;
  LAYER ME3 ;
  RECT 902.500 251.440 906.040 252.560 ;
  LAYER ME2 ;
  RECT 902.500 251.440 906.040 252.560 ;
  LAYER ME1 ;
  RECT 902.500 251.440 906.040 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 889.480 251.440 893.020 252.560 ;
  LAYER ME4 ;
  RECT 889.480 251.440 893.020 252.560 ;
  LAYER ME3 ;
  RECT 889.480 251.440 893.020 252.560 ;
  LAYER ME2 ;
  RECT 889.480 251.440 893.020 252.560 ;
  LAYER ME1 ;
  RECT 889.480 251.440 893.020 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 875.840 251.440 879.380 252.560 ;
  LAYER ME4 ;
  RECT 875.840 251.440 879.380 252.560 ;
  LAYER ME3 ;
  RECT 875.840 251.440 879.380 252.560 ;
  LAYER ME2 ;
  RECT 875.840 251.440 879.380 252.560 ;
  LAYER ME1 ;
  RECT 875.840 251.440 879.380 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 862.200 251.440 865.740 252.560 ;
  LAYER ME4 ;
  RECT 862.200 251.440 865.740 252.560 ;
  LAYER ME3 ;
  RECT 862.200 251.440 865.740 252.560 ;
  LAYER ME2 ;
  RECT 862.200 251.440 865.740 252.560 ;
  LAYER ME1 ;
  RECT 862.200 251.440 865.740 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 849.180 251.440 852.720 252.560 ;
  LAYER ME4 ;
  RECT 849.180 251.440 852.720 252.560 ;
  LAYER ME3 ;
  RECT 849.180 251.440 852.720 252.560 ;
  LAYER ME2 ;
  RECT 849.180 251.440 852.720 252.560 ;
  LAYER ME1 ;
  RECT 849.180 251.440 852.720 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 835.540 251.440 839.080 252.560 ;
  LAYER ME4 ;
  RECT 835.540 251.440 839.080 252.560 ;
  LAYER ME3 ;
  RECT 835.540 251.440 839.080 252.560 ;
  LAYER ME2 ;
  RECT 835.540 251.440 839.080 252.560 ;
  LAYER ME1 ;
  RECT 835.540 251.440 839.080 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 767.960 251.440 771.500 252.560 ;
  LAYER ME4 ;
  RECT 767.960 251.440 771.500 252.560 ;
  LAYER ME3 ;
  RECT 767.960 251.440 771.500 252.560 ;
  LAYER ME2 ;
  RECT 767.960 251.440 771.500 252.560 ;
  LAYER ME1 ;
  RECT 767.960 251.440 771.500 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 754.940 251.440 758.480 252.560 ;
  LAYER ME4 ;
  RECT 754.940 251.440 758.480 252.560 ;
  LAYER ME3 ;
  RECT 754.940 251.440 758.480 252.560 ;
  LAYER ME2 ;
  RECT 754.940 251.440 758.480 252.560 ;
  LAYER ME1 ;
  RECT 754.940 251.440 758.480 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 741.300 251.440 744.840 252.560 ;
  LAYER ME4 ;
  RECT 741.300 251.440 744.840 252.560 ;
  LAYER ME3 ;
  RECT 741.300 251.440 744.840 252.560 ;
  LAYER ME2 ;
  RECT 741.300 251.440 744.840 252.560 ;
  LAYER ME1 ;
  RECT 741.300 251.440 744.840 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 727.660 251.440 731.200 252.560 ;
  LAYER ME4 ;
  RECT 727.660 251.440 731.200 252.560 ;
  LAYER ME3 ;
  RECT 727.660 251.440 731.200 252.560 ;
  LAYER ME2 ;
  RECT 727.660 251.440 731.200 252.560 ;
  LAYER ME1 ;
  RECT 727.660 251.440 731.200 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 714.640 251.440 718.180 252.560 ;
  LAYER ME4 ;
  RECT 714.640 251.440 718.180 252.560 ;
  LAYER ME3 ;
  RECT 714.640 251.440 718.180 252.560 ;
  LAYER ME2 ;
  RECT 714.640 251.440 718.180 252.560 ;
  LAYER ME1 ;
  RECT 714.640 251.440 718.180 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 701.000 251.440 704.540 252.560 ;
  LAYER ME4 ;
  RECT 701.000 251.440 704.540 252.560 ;
  LAYER ME3 ;
  RECT 701.000 251.440 704.540 252.560 ;
  LAYER ME2 ;
  RECT 701.000 251.440 704.540 252.560 ;
  LAYER ME1 ;
  RECT 701.000 251.440 704.540 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 634.040 251.440 637.580 252.560 ;
  LAYER ME4 ;
  RECT 634.040 251.440 637.580 252.560 ;
  LAYER ME3 ;
  RECT 634.040 251.440 637.580 252.560 ;
  LAYER ME2 ;
  RECT 634.040 251.440 637.580 252.560 ;
  LAYER ME1 ;
  RECT 634.040 251.440 637.580 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 620.400 251.440 623.940 252.560 ;
  LAYER ME4 ;
  RECT 620.400 251.440 623.940 252.560 ;
  LAYER ME3 ;
  RECT 620.400 251.440 623.940 252.560 ;
  LAYER ME2 ;
  RECT 620.400 251.440 623.940 252.560 ;
  LAYER ME1 ;
  RECT 620.400 251.440 623.940 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 606.760 251.440 610.300 252.560 ;
  LAYER ME4 ;
  RECT 606.760 251.440 610.300 252.560 ;
  LAYER ME3 ;
  RECT 606.760 251.440 610.300 252.560 ;
  LAYER ME2 ;
  RECT 606.760 251.440 610.300 252.560 ;
  LAYER ME1 ;
  RECT 606.760 251.440 610.300 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 593.740 251.440 597.280 252.560 ;
  LAYER ME4 ;
  RECT 593.740 251.440 597.280 252.560 ;
  LAYER ME3 ;
  RECT 593.740 251.440 597.280 252.560 ;
  LAYER ME2 ;
  RECT 593.740 251.440 597.280 252.560 ;
  LAYER ME1 ;
  RECT 593.740 251.440 597.280 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 580.100 251.440 583.640 252.560 ;
  LAYER ME4 ;
  RECT 580.100 251.440 583.640 252.560 ;
  LAYER ME3 ;
  RECT 580.100 251.440 583.640 252.560 ;
  LAYER ME2 ;
  RECT 580.100 251.440 583.640 252.560 ;
  LAYER ME1 ;
  RECT 580.100 251.440 583.640 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 566.460 251.440 570.000 252.560 ;
  LAYER ME4 ;
  RECT 566.460 251.440 570.000 252.560 ;
  LAYER ME3 ;
  RECT 566.460 251.440 570.000 252.560 ;
  LAYER ME2 ;
  RECT 566.460 251.440 570.000 252.560 ;
  LAYER ME1 ;
  RECT 566.460 251.440 570.000 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 489.580 251.440 493.120 252.560 ;
  LAYER ME4 ;
  RECT 489.580 251.440 493.120 252.560 ;
  LAYER ME3 ;
  RECT 489.580 251.440 493.120 252.560 ;
  LAYER ME2 ;
  RECT 489.580 251.440 493.120 252.560 ;
  LAYER ME1 ;
  RECT 489.580 251.440 493.120 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 464.160 251.440 467.700 252.560 ;
  LAYER ME4 ;
  RECT 464.160 251.440 467.700 252.560 ;
  LAYER ME3 ;
  RECT 464.160 251.440 467.700 252.560 ;
  LAYER ME2 ;
  RECT 464.160 251.440 467.700 252.560 ;
  LAYER ME1 ;
  RECT 464.160 251.440 467.700 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 444.320 251.440 447.860 252.560 ;
  LAYER ME4 ;
  RECT 444.320 251.440 447.860 252.560 ;
  LAYER ME3 ;
  RECT 444.320 251.440 447.860 252.560 ;
  LAYER ME2 ;
  RECT 444.320 251.440 447.860 252.560 ;
  LAYER ME1 ;
  RECT 444.320 251.440 447.860 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 435.640 251.440 439.180 252.560 ;
  LAYER ME4 ;
  RECT 435.640 251.440 439.180 252.560 ;
  LAYER ME3 ;
  RECT 435.640 251.440 439.180 252.560 ;
  LAYER ME2 ;
  RECT 435.640 251.440 439.180 252.560 ;
  LAYER ME1 ;
  RECT 435.640 251.440 439.180 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 422.620 251.440 426.160 252.560 ;
  LAYER ME4 ;
  RECT 422.620 251.440 426.160 252.560 ;
  LAYER ME3 ;
  RECT 422.620 251.440 426.160 252.560 ;
  LAYER ME2 ;
  RECT 422.620 251.440 426.160 252.560 ;
  LAYER ME1 ;
  RECT 422.620 251.440 426.160 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 408.980 251.440 412.520 252.560 ;
  LAYER ME4 ;
  RECT 408.980 251.440 412.520 252.560 ;
  LAYER ME3 ;
  RECT 408.980 251.440 412.520 252.560 ;
  LAYER ME2 ;
  RECT 408.980 251.440 412.520 252.560 ;
  LAYER ME1 ;
  RECT 408.980 251.440 412.520 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 342.020 251.440 345.560 252.560 ;
  LAYER ME4 ;
  RECT 342.020 251.440 345.560 252.560 ;
  LAYER ME3 ;
  RECT 342.020 251.440 345.560 252.560 ;
  LAYER ME2 ;
  RECT 342.020 251.440 345.560 252.560 ;
  LAYER ME1 ;
  RECT 342.020 251.440 345.560 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 328.380 251.440 331.920 252.560 ;
  LAYER ME4 ;
  RECT 328.380 251.440 331.920 252.560 ;
  LAYER ME3 ;
  RECT 328.380 251.440 331.920 252.560 ;
  LAYER ME2 ;
  RECT 328.380 251.440 331.920 252.560 ;
  LAYER ME1 ;
  RECT 328.380 251.440 331.920 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 314.740 251.440 318.280 252.560 ;
  LAYER ME4 ;
  RECT 314.740 251.440 318.280 252.560 ;
  LAYER ME3 ;
  RECT 314.740 251.440 318.280 252.560 ;
  LAYER ME2 ;
  RECT 314.740 251.440 318.280 252.560 ;
  LAYER ME1 ;
  RECT 314.740 251.440 318.280 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 301.720 251.440 305.260 252.560 ;
  LAYER ME4 ;
  RECT 301.720 251.440 305.260 252.560 ;
  LAYER ME3 ;
  RECT 301.720 251.440 305.260 252.560 ;
  LAYER ME2 ;
  RECT 301.720 251.440 305.260 252.560 ;
  LAYER ME1 ;
  RECT 301.720 251.440 305.260 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 288.080 251.440 291.620 252.560 ;
  LAYER ME4 ;
  RECT 288.080 251.440 291.620 252.560 ;
  LAYER ME3 ;
  RECT 288.080 251.440 291.620 252.560 ;
  LAYER ME2 ;
  RECT 288.080 251.440 291.620 252.560 ;
  LAYER ME1 ;
  RECT 288.080 251.440 291.620 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 274.440 251.440 277.980 252.560 ;
  LAYER ME4 ;
  RECT 274.440 251.440 277.980 252.560 ;
  LAYER ME3 ;
  RECT 274.440 251.440 277.980 252.560 ;
  LAYER ME2 ;
  RECT 274.440 251.440 277.980 252.560 ;
  LAYER ME1 ;
  RECT 274.440 251.440 277.980 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 207.480 251.440 211.020 252.560 ;
  LAYER ME4 ;
  RECT 207.480 251.440 211.020 252.560 ;
  LAYER ME3 ;
  RECT 207.480 251.440 211.020 252.560 ;
  LAYER ME2 ;
  RECT 207.480 251.440 211.020 252.560 ;
  LAYER ME1 ;
  RECT 207.480 251.440 211.020 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 193.840 251.440 197.380 252.560 ;
  LAYER ME4 ;
  RECT 193.840 251.440 197.380 252.560 ;
  LAYER ME3 ;
  RECT 193.840 251.440 197.380 252.560 ;
  LAYER ME2 ;
  RECT 193.840 251.440 197.380 252.560 ;
  LAYER ME1 ;
  RECT 193.840 251.440 197.380 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 180.820 251.440 184.360 252.560 ;
  LAYER ME4 ;
  RECT 180.820 251.440 184.360 252.560 ;
  LAYER ME3 ;
  RECT 180.820 251.440 184.360 252.560 ;
  LAYER ME2 ;
  RECT 180.820 251.440 184.360 252.560 ;
  LAYER ME1 ;
  RECT 180.820 251.440 184.360 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 167.180 251.440 170.720 252.560 ;
  LAYER ME4 ;
  RECT 167.180 251.440 170.720 252.560 ;
  LAYER ME3 ;
  RECT 167.180 251.440 170.720 252.560 ;
  LAYER ME2 ;
  RECT 167.180 251.440 170.720 252.560 ;
  LAYER ME1 ;
  RECT 167.180 251.440 170.720 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 153.540 251.440 157.080 252.560 ;
  LAYER ME4 ;
  RECT 153.540 251.440 157.080 252.560 ;
  LAYER ME3 ;
  RECT 153.540 251.440 157.080 252.560 ;
  LAYER ME2 ;
  RECT 153.540 251.440 157.080 252.560 ;
  LAYER ME1 ;
  RECT 153.540 251.440 157.080 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 140.520 251.440 144.060 252.560 ;
  LAYER ME4 ;
  RECT 140.520 251.440 144.060 252.560 ;
  LAYER ME3 ;
  RECT 140.520 251.440 144.060 252.560 ;
  LAYER ME2 ;
  RECT 140.520 251.440 144.060 252.560 ;
  LAYER ME1 ;
  RECT 140.520 251.440 144.060 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 72.940 251.440 76.480 252.560 ;
  LAYER ME4 ;
  RECT 72.940 251.440 76.480 252.560 ;
  LAYER ME3 ;
  RECT 72.940 251.440 76.480 252.560 ;
  LAYER ME2 ;
  RECT 72.940 251.440 76.480 252.560 ;
  LAYER ME1 ;
  RECT 72.940 251.440 76.480 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 59.300 251.440 62.840 252.560 ;
  LAYER ME4 ;
  RECT 59.300 251.440 62.840 252.560 ;
  LAYER ME3 ;
  RECT 59.300 251.440 62.840 252.560 ;
  LAYER ME2 ;
  RECT 59.300 251.440 62.840 252.560 ;
  LAYER ME1 ;
  RECT 59.300 251.440 62.840 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 46.280 251.440 49.820 252.560 ;
  LAYER ME4 ;
  RECT 46.280 251.440 49.820 252.560 ;
  LAYER ME3 ;
  RECT 46.280 251.440 49.820 252.560 ;
  LAYER ME2 ;
  RECT 46.280 251.440 49.820 252.560 ;
  LAYER ME1 ;
  RECT 46.280 251.440 49.820 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 32.640 251.440 36.180 252.560 ;
  LAYER ME4 ;
  RECT 32.640 251.440 36.180 252.560 ;
  LAYER ME3 ;
  RECT 32.640 251.440 36.180 252.560 ;
  LAYER ME2 ;
  RECT 32.640 251.440 36.180 252.560 ;
  LAYER ME1 ;
  RECT 32.640 251.440 36.180 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 19.000 251.440 22.540 252.560 ;
  LAYER ME4 ;
  RECT 19.000 251.440 22.540 252.560 ;
  LAYER ME3 ;
  RECT 19.000 251.440 22.540 252.560 ;
  LAYER ME2 ;
  RECT 19.000 251.440 22.540 252.560 ;
  LAYER ME1 ;
  RECT 19.000 251.440 22.540 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 7.220 251.440 10.760 252.560 ;
  LAYER ME4 ;
  RECT 7.220 251.440 10.760 252.560 ;
  LAYER ME3 ;
  RECT 7.220 251.440 10.760 252.560 ;
  LAYER ME2 ;
  RECT 7.220 251.440 10.760 252.560 ;
  LAYER ME1 ;
  RECT 7.220 251.440 10.760 252.560 ;
 END
 PORT
  LAYER ME5 ;
  RECT 902.500 0.000 906.040 1.120 ;
  LAYER ME4 ;
  RECT 902.500 0.000 906.040 1.120 ;
  LAYER ME3 ;
  RECT 902.500 0.000 906.040 1.120 ;
  LAYER ME2 ;
  RECT 902.500 0.000 906.040 1.120 ;
  LAYER ME1 ;
  RECT 902.500 0.000 906.040 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 889.480 0.000 893.020 1.120 ;
  LAYER ME4 ;
  RECT 889.480 0.000 893.020 1.120 ;
  LAYER ME3 ;
  RECT 889.480 0.000 893.020 1.120 ;
  LAYER ME2 ;
  RECT 889.480 0.000 893.020 1.120 ;
  LAYER ME1 ;
  RECT 889.480 0.000 893.020 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 875.840 0.000 879.380 1.120 ;
  LAYER ME4 ;
  RECT 875.840 0.000 879.380 1.120 ;
  LAYER ME3 ;
  RECT 875.840 0.000 879.380 1.120 ;
  LAYER ME2 ;
  RECT 875.840 0.000 879.380 1.120 ;
  LAYER ME1 ;
  RECT 875.840 0.000 879.380 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 862.200 0.000 865.740 1.120 ;
  LAYER ME4 ;
  RECT 862.200 0.000 865.740 1.120 ;
  LAYER ME3 ;
  RECT 862.200 0.000 865.740 1.120 ;
  LAYER ME2 ;
  RECT 862.200 0.000 865.740 1.120 ;
  LAYER ME1 ;
  RECT 862.200 0.000 865.740 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 849.180 0.000 852.720 1.120 ;
  LAYER ME4 ;
  RECT 849.180 0.000 852.720 1.120 ;
  LAYER ME3 ;
  RECT 849.180 0.000 852.720 1.120 ;
  LAYER ME2 ;
  RECT 849.180 0.000 852.720 1.120 ;
  LAYER ME1 ;
  RECT 849.180 0.000 852.720 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 835.540 0.000 839.080 1.120 ;
  LAYER ME4 ;
  RECT 835.540 0.000 839.080 1.120 ;
  LAYER ME3 ;
  RECT 835.540 0.000 839.080 1.120 ;
  LAYER ME2 ;
  RECT 835.540 0.000 839.080 1.120 ;
  LAYER ME1 ;
  RECT 835.540 0.000 839.080 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 767.960 0.000 771.500 1.120 ;
  LAYER ME4 ;
  RECT 767.960 0.000 771.500 1.120 ;
  LAYER ME3 ;
  RECT 767.960 0.000 771.500 1.120 ;
  LAYER ME2 ;
  RECT 767.960 0.000 771.500 1.120 ;
  LAYER ME1 ;
  RECT 767.960 0.000 771.500 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 754.940 0.000 758.480 1.120 ;
  LAYER ME4 ;
  RECT 754.940 0.000 758.480 1.120 ;
  LAYER ME3 ;
  RECT 754.940 0.000 758.480 1.120 ;
  LAYER ME2 ;
  RECT 754.940 0.000 758.480 1.120 ;
  LAYER ME1 ;
  RECT 754.940 0.000 758.480 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 741.300 0.000 744.840 1.120 ;
  LAYER ME4 ;
  RECT 741.300 0.000 744.840 1.120 ;
  LAYER ME3 ;
  RECT 741.300 0.000 744.840 1.120 ;
  LAYER ME2 ;
  RECT 741.300 0.000 744.840 1.120 ;
  LAYER ME1 ;
  RECT 741.300 0.000 744.840 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 727.660 0.000 731.200 1.120 ;
  LAYER ME4 ;
  RECT 727.660 0.000 731.200 1.120 ;
  LAYER ME3 ;
  RECT 727.660 0.000 731.200 1.120 ;
  LAYER ME2 ;
  RECT 727.660 0.000 731.200 1.120 ;
  LAYER ME1 ;
  RECT 727.660 0.000 731.200 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 714.640 0.000 718.180 1.120 ;
  LAYER ME4 ;
  RECT 714.640 0.000 718.180 1.120 ;
  LAYER ME3 ;
  RECT 714.640 0.000 718.180 1.120 ;
  LAYER ME2 ;
  RECT 714.640 0.000 718.180 1.120 ;
  LAYER ME1 ;
  RECT 714.640 0.000 718.180 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 701.000 0.000 704.540 1.120 ;
  LAYER ME4 ;
  RECT 701.000 0.000 704.540 1.120 ;
  LAYER ME3 ;
  RECT 701.000 0.000 704.540 1.120 ;
  LAYER ME2 ;
  RECT 701.000 0.000 704.540 1.120 ;
  LAYER ME1 ;
  RECT 701.000 0.000 704.540 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 634.040 0.000 637.580 1.120 ;
  LAYER ME4 ;
  RECT 634.040 0.000 637.580 1.120 ;
  LAYER ME3 ;
  RECT 634.040 0.000 637.580 1.120 ;
  LAYER ME2 ;
  RECT 634.040 0.000 637.580 1.120 ;
  LAYER ME1 ;
  RECT 634.040 0.000 637.580 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 620.400 0.000 623.940 1.120 ;
  LAYER ME4 ;
  RECT 620.400 0.000 623.940 1.120 ;
  LAYER ME3 ;
  RECT 620.400 0.000 623.940 1.120 ;
  LAYER ME2 ;
  RECT 620.400 0.000 623.940 1.120 ;
  LAYER ME1 ;
  RECT 620.400 0.000 623.940 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 606.760 0.000 610.300 1.120 ;
  LAYER ME4 ;
  RECT 606.760 0.000 610.300 1.120 ;
  LAYER ME3 ;
  RECT 606.760 0.000 610.300 1.120 ;
  LAYER ME2 ;
  RECT 606.760 0.000 610.300 1.120 ;
  LAYER ME1 ;
  RECT 606.760 0.000 610.300 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 593.740 0.000 597.280 1.120 ;
  LAYER ME4 ;
  RECT 593.740 0.000 597.280 1.120 ;
  LAYER ME3 ;
  RECT 593.740 0.000 597.280 1.120 ;
  LAYER ME2 ;
  RECT 593.740 0.000 597.280 1.120 ;
  LAYER ME1 ;
  RECT 593.740 0.000 597.280 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 580.100 0.000 583.640 1.120 ;
  LAYER ME4 ;
  RECT 580.100 0.000 583.640 1.120 ;
  LAYER ME3 ;
  RECT 580.100 0.000 583.640 1.120 ;
  LAYER ME2 ;
  RECT 580.100 0.000 583.640 1.120 ;
  LAYER ME1 ;
  RECT 580.100 0.000 583.640 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 566.460 0.000 570.000 1.120 ;
  LAYER ME4 ;
  RECT 566.460 0.000 570.000 1.120 ;
  LAYER ME3 ;
  RECT 566.460 0.000 570.000 1.120 ;
  LAYER ME2 ;
  RECT 566.460 0.000 570.000 1.120 ;
  LAYER ME1 ;
  RECT 566.460 0.000 570.000 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 489.580 0.000 493.120 1.120 ;
  LAYER ME4 ;
  RECT 489.580 0.000 493.120 1.120 ;
  LAYER ME3 ;
  RECT 489.580 0.000 493.120 1.120 ;
  LAYER ME2 ;
  RECT 489.580 0.000 493.120 1.120 ;
  LAYER ME1 ;
  RECT 489.580 0.000 493.120 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 464.160 0.000 467.700 1.120 ;
  LAYER ME4 ;
  RECT 464.160 0.000 467.700 1.120 ;
  LAYER ME3 ;
  RECT 464.160 0.000 467.700 1.120 ;
  LAYER ME2 ;
  RECT 464.160 0.000 467.700 1.120 ;
  LAYER ME1 ;
  RECT 464.160 0.000 467.700 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 444.320 0.000 447.860 1.120 ;
  LAYER ME4 ;
  RECT 444.320 0.000 447.860 1.120 ;
  LAYER ME3 ;
  RECT 444.320 0.000 447.860 1.120 ;
  LAYER ME2 ;
  RECT 444.320 0.000 447.860 1.120 ;
  LAYER ME1 ;
  RECT 444.320 0.000 447.860 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 435.640 0.000 439.180 1.120 ;
  LAYER ME4 ;
  RECT 435.640 0.000 439.180 1.120 ;
  LAYER ME3 ;
  RECT 435.640 0.000 439.180 1.120 ;
  LAYER ME2 ;
  RECT 435.640 0.000 439.180 1.120 ;
  LAYER ME1 ;
  RECT 435.640 0.000 439.180 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 422.620 0.000 426.160 1.120 ;
  LAYER ME4 ;
  RECT 422.620 0.000 426.160 1.120 ;
  LAYER ME3 ;
  RECT 422.620 0.000 426.160 1.120 ;
  LAYER ME2 ;
  RECT 422.620 0.000 426.160 1.120 ;
  LAYER ME1 ;
  RECT 422.620 0.000 426.160 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 408.980 0.000 412.520 1.120 ;
  LAYER ME4 ;
  RECT 408.980 0.000 412.520 1.120 ;
  LAYER ME3 ;
  RECT 408.980 0.000 412.520 1.120 ;
  LAYER ME2 ;
  RECT 408.980 0.000 412.520 1.120 ;
  LAYER ME1 ;
  RECT 408.980 0.000 412.520 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 342.020 0.000 345.560 1.120 ;
  LAYER ME4 ;
  RECT 342.020 0.000 345.560 1.120 ;
  LAYER ME3 ;
  RECT 342.020 0.000 345.560 1.120 ;
  LAYER ME2 ;
  RECT 342.020 0.000 345.560 1.120 ;
  LAYER ME1 ;
  RECT 342.020 0.000 345.560 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 328.380 0.000 331.920 1.120 ;
  LAYER ME4 ;
  RECT 328.380 0.000 331.920 1.120 ;
  LAYER ME3 ;
  RECT 328.380 0.000 331.920 1.120 ;
  LAYER ME2 ;
  RECT 328.380 0.000 331.920 1.120 ;
  LAYER ME1 ;
  RECT 328.380 0.000 331.920 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 314.740 0.000 318.280 1.120 ;
  LAYER ME4 ;
  RECT 314.740 0.000 318.280 1.120 ;
  LAYER ME3 ;
  RECT 314.740 0.000 318.280 1.120 ;
  LAYER ME2 ;
  RECT 314.740 0.000 318.280 1.120 ;
  LAYER ME1 ;
  RECT 314.740 0.000 318.280 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 301.720 0.000 305.260 1.120 ;
  LAYER ME4 ;
  RECT 301.720 0.000 305.260 1.120 ;
  LAYER ME3 ;
  RECT 301.720 0.000 305.260 1.120 ;
  LAYER ME2 ;
  RECT 301.720 0.000 305.260 1.120 ;
  LAYER ME1 ;
  RECT 301.720 0.000 305.260 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 288.080 0.000 291.620 1.120 ;
  LAYER ME4 ;
  RECT 288.080 0.000 291.620 1.120 ;
  LAYER ME3 ;
  RECT 288.080 0.000 291.620 1.120 ;
  LAYER ME2 ;
  RECT 288.080 0.000 291.620 1.120 ;
  LAYER ME1 ;
  RECT 288.080 0.000 291.620 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 274.440 0.000 277.980 1.120 ;
  LAYER ME4 ;
  RECT 274.440 0.000 277.980 1.120 ;
  LAYER ME3 ;
  RECT 274.440 0.000 277.980 1.120 ;
  LAYER ME2 ;
  RECT 274.440 0.000 277.980 1.120 ;
  LAYER ME1 ;
  RECT 274.440 0.000 277.980 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 207.480 0.000 211.020 1.120 ;
  LAYER ME4 ;
  RECT 207.480 0.000 211.020 1.120 ;
  LAYER ME3 ;
  RECT 207.480 0.000 211.020 1.120 ;
  LAYER ME2 ;
  RECT 207.480 0.000 211.020 1.120 ;
  LAYER ME1 ;
  RECT 207.480 0.000 211.020 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 193.840 0.000 197.380 1.120 ;
  LAYER ME4 ;
  RECT 193.840 0.000 197.380 1.120 ;
  LAYER ME3 ;
  RECT 193.840 0.000 197.380 1.120 ;
  LAYER ME2 ;
  RECT 193.840 0.000 197.380 1.120 ;
  LAYER ME1 ;
  RECT 193.840 0.000 197.380 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 180.820 0.000 184.360 1.120 ;
  LAYER ME4 ;
  RECT 180.820 0.000 184.360 1.120 ;
  LAYER ME3 ;
  RECT 180.820 0.000 184.360 1.120 ;
  LAYER ME2 ;
  RECT 180.820 0.000 184.360 1.120 ;
  LAYER ME1 ;
  RECT 180.820 0.000 184.360 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 167.180 0.000 170.720 1.120 ;
  LAYER ME4 ;
  RECT 167.180 0.000 170.720 1.120 ;
  LAYER ME3 ;
  RECT 167.180 0.000 170.720 1.120 ;
  LAYER ME2 ;
  RECT 167.180 0.000 170.720 1.120 ;
  LAYER ME1 ;
  RECT 167.180 0.000 170.720 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 153.540 0.000 157.080 1.120 ;
  LAYER ME4 ;
  RECT 153.540 0.000 157.080 1.120 ;
  LAYER ME3 ;
  RECT 153.540 0.000 157.080 1.120 ;
  LAYER ME2 ;
  RECT 153.540 0.000 157.080 1.120 ;
  LAYER ME1 ;
  RECT 153.540 0.000 157.080 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 140.520 0.000 144.060 1.120 ;
  LAYER ME4 ;
  RECT 140.520 0.000 144.060 1.120 ;
  LAYER ME3 ;
  RECT 140.520 0.000 144.060 1.120 ;
  LAYER ME2 ;
  RECT 140.520 0.000 144.060 1.120 ;
  LAYER ME1 ;
  RECT 140.520 0.000 144.060 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 72.940 0.000 76.480 1.120 ;
  LAYER ME4 ;
  RECT 72.940 0.000 76.480 1.120 ;
  LAYER ME3 ;
  RECT 72.940 0.000 76.480 1.120 ;
  LAYER ME2 ;
  RECT 72.940 0.000 76.480 1.120 ;
  LAYER ME1 ;
  RECT 72.940 0.000 76.480 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 59.300 0.000 62.840 1.120 ;
  LAYER ME4 ;
  RECT 59.300 0.000 62.840 1.120 ;
  LAYER ME3 ;
  RECT 59.300 0.000 62.840 1.120 ;
  LAYER ME2 ;
  RECT 59.300 0.000 62.840 1.120 ;
  LAYER ME1 ;
  RECT 59.300 0.000 62.840 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 46.280 0.000 49.820 1.120 ;
  LAYER ME4 ;
  RECT 46.280 0.000 49.820 1.120 ;
  LAYER ME3 ;
  RECT 46.280 0.000 49.820 1.120 ;
  LAYER ME2 ;
  RECT 46.280 0.000 49.820 1.120 ;
  LAYER ME1 ;
  RECT 46.280 0.000 49.820 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 32.640 0.000 36.180 1.120 ;
  LAYER ME4 ;
  RECT 32.640 0.000 36.180 1.120 ;
  LAYER ME3 ;
  RECT 32.640 0.000 36.180 1.120 ;
  LAYER ME2 ;
  RECT 32.640 0.000 36.180 1.120 ;
  LAYER ME1 ;
  RECT 32.640 0.000 36.180 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 19.000 0.000 22.540 1.120 ;
  LAYER ME4 ;
  RECT 19.000 0.000 22.540 1.120 ;
  LAYER ME3 ;
  RECT 19.000 0.000 22.540 1.120 ;
  LAYER ME2 ;
  RECT 19.000 0.000 22.540 1.120 ;
  LAYER ME1 ;
  RECT 19.000 0.000 22.540 1.120 ;
 END
 PORT
  LAYER ME5 ;
  RECT 7.220 0.000 10.760 1.120 ;
  LAYER ME4 ;
  RECT 7.220 0.000 10.760 1.120 ;
  LAYER ME3 ;
  RECT 7.220 0.000 10.760 1.120 ;
  LAYER ME2 ;
  RECT 7.220 0.000 10.760 1.120 ;
  LAYER ME1 ;
  RECT 7.220 0.000 10.760 1.120 ;
 END
END VCC
PIN DIB31
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER ME5 ;
  RECT 949.900 251.440 951.020 252.560 ;
  LAYER ME4 ;
  RECT 949.900 251.440 951.020 252.560 ;
  LAYER ME3 ;
  RECT 949.900 251.440 951.020 252.560 ;
  LAYER ME2 ;
  RECT 949.900 251.440 951.020 252.560 ;
  LAYER ME1 ;
  RECT 949.900 251.440 951.020 252.560 ;
 END
END DIB31
PIN DOB31
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME5 ;
  RECT 936.260 251.440 937.380 252.560 ;
  LAYER ME4 ;
  RECT 936.260 251.440 937.380 252.560 ;
  LAYER ME3 ;
  RECT 936.260 251.440 937.380 252.560 ;
  LAYER ME2 ;
  RECT 936.260 251.440 937.380 252.560 ;
  LAYER ME1 ;
  RECT 936.260 251.440 937.380 252.560 ;
 END
END DOB31
PIN DIB30
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER ME5 ;
  RECT 923.240 251.440 924.360 252.560 ;
  LAYER ME4 ;
  RECT 923.240 251.440 924.360 252.560 ;
  LAYER ME3 ;
  RECT 923.240 251.440 924.360 252.560 ;
  LAYER ME2 ;
  RECT 923.240 251.440 924.360 252.560 ;
  LAYER ME1 ;
  RECT 923.240 251.440 924.360 252.560 ;
 END
END DIB30
PIN DOB30
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME5 ;
  RECT 909.600 251.440 910.720 252.560 ;
  LAYER ME4 ;
  RECT 909.600 251.440 910.720 252.560 ;
  LAYER ME3 ;
  RECT 909.600 251.440 910.720 252.560 ;
  LAYER ME2 ;
  RECT 909.600 251.440 910.720 252.560 ;
  LAYER ME1 ;
  RECT 909.600 251.440 910.720 252.560 ;
 END
END DOB30
PIN DIB29
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER ME5 ;
  RECT 895.960 251.440 897.080 252.560 ;
  LAYER ME4 ;
  RECT 895.960 251.440 897.080 252.560 ;
  LAYER ME3 ;
  RECT 895.960 251.440 897.080 252.560 ;
  LAYER ME2 ;
  RECT 895.960 251.440 897.080 252.560 ;
  LAYER ME1 ;
  RECT 895.960 251.440 897.080 252.560 ;
 END
END DIB29
PIN DOB29
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME5 ;
  RECT 882.940 251.440 884.060 252.560 ;
  LAYER ME4 ;
  RECT 882.940 251.440 884.060 252.560 ;
  LAYER ME3 ;
  RECT 882.940 251.440 884.060 252.560 ;
  LAYER ME2 ;
  RECT 882.940 251.440 884.060 252.560 ;
  LAYER ME1 ;
  RECT 882.940 251.440 884.060 252.560 ;
 END
END DOB29
PIN DIB28
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER ME5 ;
  RECT 869.300 251.440 870.420 252.560 ;
  LAYER ME4 ;
  RECT 869.300 251.440 870.420 252.560 ;
  LAYER ME3 ;
  RECT 869.300 251.440 870.420 252.560 ;
  LAYER ME2 ;
  RECT 869.300 251.440 870.420 252.560 ;
  LAYER ME1 ;
  RECT 869.300 251.440 870.420 252.560 ;
 END
END DIB28
PIN DOB28
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME5 ;
  RECT 855.660 251.440 856.780 252.560 ;
  LAYER ME4 ;
  RECT 855.660 251.440 856.780 252.560 ;
  LAYER ME3 ;
  RECT 855.660 251.440 856.780 252.560 ;
  LAYER ME2 ;
  RECT 855.660 251.440 856.780 252.560 ;
  LAYER ME1 ;
  RECT 855.660 251.440 856.780 252.560 ;
 END
END DOB28
PIN DIB27
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER ME5 ;
  RECT 842.640 251.440 843.760 252.560 ;
  LAYER ME4 ;
  RECT 842.640 251.440 843.760 252.560 ;
  LAYER ME3 ;
  RECT 842.640 251.440 843.760 252.560 ;
  LAYER ME2 ;
  RECT 842.640 251.440 843.760 252.560 ;
  LAYER ME1 ;
  RECT 842.640 251.440 843.760 252.560 ;
 END
END DIB27
PIN DOB27
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME5 ;
  RECT 829.000 251.440 830.120 252.560 ;
  LAYER ME4 ;
  RECT 829.000 251.440 830.120 252.560 ;
  LAYER ME3 ;
  RECT 829.000 251.440 830.120 252.560 ;
  LAYER ME2 ;
  RECT 829.000 251.440 830.120 252.560 ;
  LAYER ME1 ;
  RECT 829.000 251.440 830.120 252.560 ;
 END
END DOB27
PIN DIB26
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER ME5 ;
  RECT 815.360 251.440 816.480 252.560 ;
  LAYER ME4 ;
  RECT 815.360 251.440 816.480 252.560 ;
  LAYER ME3 ;
  RECT 815.360 251.440 816.480 252.560 ;
  LAYER ME2 ;
  RECT 815.360 251.440 816.480 252.560 ;
  LAYER ME1 ;
  RECT 815.360 251.440 816.480 252.560 ;
 END
END DIB26
PIN DOB26
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME5 ;
  RECT 802.340 251.440 803.460 252.560 ;
  LAYER ME4 ;
  RECT 802.340 251.440 803.460 252.560 ;
  LAYER ME3 ;
  RECT 802.340 251.440 803.460 252.560 ;
  LAYER ME2 ;
  RECT 802.340 251.440 803.460 252.560 ;
  LAYER ME1 ;
  RECT 802.340 251.440 803.460 252.560 ;
 END
END DOB26
PIN DIB25
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER ME5 ;
  RECT 788.700 251.440 789.820 252.560 ;
  LAYER ME4 ;
  RECT 788.700 251.440 789.820 252.560 ;
  LAYER ME3 ;
  RECT 788.700 251.440 789.820 252.560 ;
  LAYER ME2 ;
  RECT 788.700 251.440 789.820 252.560 ;
  LAYER ME1 ;
  RECT 788.700 251.440 789.820 252.560 ;
 END
END DIB25
PIN DOB25
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME5 ;
  RECT 775.060 251.440 776.180 252.560 ;
  LAYER ME4 ;
  RECT 775.060 251.440 776.180 252.560 ;
  LAYER ME3 ;
  RECT 775.060 251.440 776.180 252.560 ;
  LAYER ME2 ;
  RECT 775.060 251.440 776.180 252.560 ;
  LAYER ME1 ;
  RECT 775.060 251.440 776.180 252.560 ;
 END
END DOB25
PIN DIB24
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER ME5 ;
  RECT 761.420 251.440 762.540 252.560 ;
  LAYER ME4 ;
  RECT 761.420 251.440 762.540 252.560 ;
  LAYER ME3 ;
  RECT 761.420 251.440 762.540 252.560 ;
  LAYER ME2 ;
  RECT 761.420 251.440 762.540 252.560 ;
  LAYER ME1 ;
  RECT 761.420 251.440 762.540 252.560 ;
 END
END DIB24
PIN DOB24
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME5 ;
  RECT 748.400 251.440 749.520 252.560 ;
  LAYER ME4 ;
  RECT 748.400 251.440 749.520 252.560 ;
  LAYER ME3 ;
  RECT 748.400 251.440 749.520 252.560 ;
  LAYER ME2 ;
  RECT 748.400 251.440 749.520 252.560 ;
  LAYER ME1 ;
  RECT 748.400 251.440 749.520 252.560 ;
 END
END DOB24
PIN DIB23
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER ME5 ;
  RECT 734.760 251.440 735.880 252.560 ;
  LAYER ME4 ;
  RECT 734.760 251.440 735.880 252.560 ;
  LAYER ME3 ;
  RECT 734.760 251.440 735.880 252.560 ;
  LAYER ME2 ;
  RECT 734.760 251.440 735.880 252.560 ;
  LAYER ME1 ;
  RECT 734.760 251.440 735.880 252.560 ;
 END
END DIB23
PIN DOB23
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME5 ;
  RECT 721.120 251.440 722.240 252.560 ;
  LAYER ME4 ;
  RECT 721.120 251.440 722.240 252.560 ;
  LAYER ME3 ;
  RECT 721.120 251.440 722.240 252.560 ;
  LAYER ME2 ;
  RECT 721.120 251.440 722.240 252.560 ;
  LAYER ME1 ;
  RECT 721.120 251.440 722.240 252.560 ;
 END
END DOB23
PIN DIB22
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER ME5 ;
  RECT 708.100 251.440 709.220 252.560 ;
  LAYER ME4 ;
  RECT 708.100 251.440 709.220 252.560 ;
  LAYER ME3 ;
  RECT 708.100 251.440 709.220 252.560 ;
  LAYER ME2 ;
  RECT 708.100 251.440 709.220 252.560 ;
  LAYER ME1 ;
  RECT 708.100 251.440 709.220 252.560 ;
 END
END DIB22
PIN DOB22
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME5 ;
  RECT 694.460 251.440 695.580 252.560 ;
  LAYER ME4 ;
  RECT 694.460 251.440 695.580 252.560 ;
  LAYER ME3 ;
  RECT 694.460 251.440 695.580 252.560 ;
  LAYER ME2 ;
  RECT 694.460 251.440 695.580 252.560 ;
  LAYER ME1 ;
  RECT 694.460 251.440 695.580 252.560 ;
 END
END DOB22
PIN DIB21
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER ME5 ;
  RECT 680.820 251.440 681.940 252.560 ;
  LAYER ME4 ;
  RECT 680.820 251.440 681.940 252.560 ;
  LAYER ME3 ;
  RECT 680.820 251.440 681.940 252.560 ;
  LAYER ME2 ;
  RECT 680.820 251.440 681.940 252.560 ;
  LAYER ME1 ;
  RECT 680.820 251.440 681.940 252.560 ;
 END
END DIB21
PIN DOB21
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME5 ;
  RECT 667.800 251.440 668.920 252.560 ;
  LAYER ME4 ;
  RECT 667.800 251.440 668.920 252.560 ;
  LAYER ME3 ;
  RECT 667.800 251.440 668.920 252.560 ;
  LAYER ME2 ;
  RECT 667.800 251.440 668.920 252.560 ;
  LAYER ME1 ;
  RECT 667.800 251.440 668.920 252.560 ;
 END
END DOB21
PIN DIB20
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER ME5 ;
  RECT 654.160 251.440 655.280 252.560 ;
  LAYER ME4 ;
  RECT 654.160 251.440 655.280 252.560 ;
  LAYER ME3 ;
  RECT 654.160 251.440 655.280 252.560 ;
  LAYER ME2 ;
  RECT 654.160 251.440 655.280 252.560 ;
  LAYER ME1 ;
  RECT 654.160 251.440 655.280 252.560 ;
 END
END DIB20
PIN DOB20
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME5 ;
  RECT 640.520 251.440 641.640 252.560 ;
  LAYER ME4 ;
  RECT 640.520 251.440 641.640 252.560 ;
  LAYER ME3 ;
  RECT 640.520 251.440 641.640 252.560 ;
  LAYER ME2 ;
  RECT 640.520 251.440 641.640 252.560 ;
  LAYER ME1 ;
  RECT 640.520 251.440 641.640 252.560 ;
 END
END DOB20
PIN DIB19
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER ME5 ;
  RECT 627.500 251.440 628.620 252.560 ;
  LAYER ME4 ;
  RECT 627.500 251.440 628.620 252.560 ;
  LAYER ME3 ;
  RECT 627.500 251.440 628.620 252.560 ;
  LAYER ME2 ;
  RECT 627.500 251.440 628.620 252.560 ;
  LAYER ME1 ;
  RECT 627.500 251.440 628.620 252.560 ;
 END
END DIB19
PIN DOB19
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME5 ;
  RECT 613.860 251.440 614.980 252.560 ;
  LAYER ME4 ;
  RECT 613.860 251.440 614.980 252.560 ;
  LAYER ME3 ;
  RECT 613.860 251.440 614.980 252.560 ;
  LAYER ME2 ;
  RECT 613.860 251.440 614.980 252.560 ;
  LAYER ME1 ;
  RECT 613.860 251.440 614.980 252.560 ;
 END
END DOB19
PIN DIB18
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER ME5 ;
  RECT 600.220 251.440 601.340 252.560 ;
  LAYER ME4 ;
  RECT 600.220 251.440 601.340 252.560 ;
  LAYER ME3 ;
  RECT 600.220 251.440 601.340 252.560 ;
  LAYER ME2 ;
  RECT 600.220 251.440 601.340 252.560 ;
  LAYER ME1 ;
  RECT 600.220 251.440 601.340 252.560 ;
 END
END DIB18
PIN DOB18
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME5 ;
  RECT 587.200 251.440 588.320 252.560 ;
  LAYER ME4 ;
  RECT 587.200 251.440 588.320 252.560 ;
  LAYER ME3 ;
  RECT 587.200 251.440 588.320 252.560 ;
  LAYER ME2 ;
  RECT 587.200 251.440 588.320 252.560 ;
  LAYER ME1 ;
  RECT 587.200 251.440 588.320 252.560 ;
 END
END DOB18
PIN DIB17
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER ME5 ;
  RECT 573.560 251.440 574.680 252.560 ;
  LAYER ME4 ;
  RECT 573.560 251.440 574.680 252.560 ;
  LAYER ME3 ;
  RECT 573.560 251.440 574.680 252.560 ;
  LAYER ME2 ;
  RECT 573.560 251.440 574.680 252.560 ;
  LAYER ME1 ;
  RECT 573.560 251.440 574.680 252.560 ;
 END
END DIB17
PIN DOB17
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME5 ;
  RECT 559.920 251.440 561.040 252.560 ;
  LAYER ME4 ;
  RECT 559.920 251.440 561.040 252.560 ;
  LAYER ME3 ;
  RECT 559.920 251.440 561.040 252.560 ;
  LAYER ME2 ;
  RECT 559.920 251.440 561.040 252.560 ;
  LAYER ME1 ;
  RECT 559.920 251.440 561.040 252.560 ;
 END
END DOB17
PIN DIB16
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER ME5 ;
  RECT 546.900 251.440 548.020 252.560 ;
  LAYER ME4 ;
  RECT 546.900 251.440 548.020 252.560 ;
  LAYER ME3 ;
  RECT 546.900 251.440 548.020 252.560 ;
  LAYER ME2 ;
  RECT 546.900 251.440 548.020 252.560 ;
  LAYER ME1 ;
  RECT 546.900 251.440 548.020 252.560 ;
 END
END DIB16
PIN DOB16
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME5 ;
  RECT 533.260 251.440 534.380 252.560 ;
  LAYER ME4 ;
  RECT 533.260 251.440 534.380 252.560 ;
  LAYER ME3 ;
  RECT 533.260 251.440 534.380 252.560 ;
  LAYER ME2 ;
  RECT 533.260 251.440 534.380 252.560 ;
  LAYER ME1 ;
  RECT 533.260 251.440 534.380 252.560 ;
 END
END DOB16
PIN CKB
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER ME5 ;
  RECT 511.560 251.440 512.680 252.560 ;
  LAYER ME4 ;
  RECT 511.560 251.440 512.680 252.560 ;
  LAYER ME3 ;
  RECT 511.560 251.440 512.680 252.560 ;
  LAYER ME2 ;
  RECT 511.560 251.440 512.680 252.560 ;
  LAYER ME1 ;
  RECT 511.560 251.440 512.680 252.560 ;
 END
END CKB
PIN CSB
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER ME5 ;
  RECT 509.080 251.440 510.200 252.560 ;
  LAYER ME4 ;
  RECT 509.080 251.440 510.200 252.560 ;
  LAYER ME3 ;
  RECT 509.080 251.440 510.200 252.560 ;
  LAYER ME2 ;
  RECT 509.080 251.440 510.200 252.560 ;
  LAYER ME1 ;
  RECT 509.080 251.440 510.200 252.560 ;
 END
END CSB
PIN WEBN
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER ME5 ;
  RECT 507.220 251.440 508.340 252.560 ;
  LAYER ME4 ;
  RECT 507.220 251.440 508.340 252.560 ;
  LAYER ME3 ;
  RECT 507.220 251.440 508.340 252.560 ;
  LAYER ME2 ;
  RECT 507.220 251.440 508.340 252.560 ;
  LAYER ME1 ;
  RECT 507.220 251.440 508.340 252.560 ;
 END
END WEBN
PIN B2
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER ME5 ;
  RECT 503.500 251.440 504.620 252.560 ;
  LAYER ME4 ;
  RECT 503.500 251.440 504.620 252.560 ;
  LAYER ME3 ;
  RECT 503.500 251.440 504.620 252.560 ;
  LAYER ME2 ;
  RECT 503.500 251.440 504.620 252.560 ;
  LAYER ME1 ;
  RECT 503.500 251.440 504.620 252.560 ;
 END
END B2
PIN OEB
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER ME5 ;
  RECT 499.780 251.440 500.900 252.560 ;
  LAYER ME4 ;
  RECT 499.780 251.440 500.900 252.560 ;
  LAYER ME3 ;
  RECT 499.780 251.440 500.900 252.560 ;
  LAYER ME2 ;
  RECT 499.780 251.440 500.900 252.560 ;
  LAYER ME1 ;
  RECT 499.780 251.440 500.900 252.560 ;
 END
END OEB
PIN B1
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER ME5 ;
  RECT 497.920 251.440 499.040 252.560 ;
  LAYER ME4 ;
  RECT 497.920 251.440 499.040 252.560 ;
  LAYER ME3 ;
  RECT 497.920 251.440 499.040 252.560 ;
  LAYER ME2 ;
  RECT 497.920 251.440 499.040 252.560 ;
  LAYER ME1 ;
  RECT 497.920 251.440 499.040 252.560 ;
 END
END B1
PIN B0
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER ME5 ;
  RECT 496.060 251.440 497.180 252.560 ;
  LAYER ME4 ;
  RECT 496.060 251.440 497.180 252.560 ;
  LAYER ME3 ;
  RECT 496.060 251.440 497.180 252.560 ;
  LAYER ME2 ;
  RECT 496.060 251.440 497.180 252.560 ;
  LAYER ME1 ;
  RECT 496.060 251.440 497.180 252.560 ;
 END
END B0
PIN B5
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER ME5 ;
  RECT 487.380 251.440 488.500 252.560 ;
  LAYER ME4 ;
  RECT 487.380 251.440 488.500 252.560 ;
  LAYER ME3 ;
  RECT 487.380 251.440 488.500 252.560 ;
  LAYER ME2 ;
  RECT 487.380 251.440 488.500 252.560 ;
  LAYER ME1 ;
  RECT 487.380 251.440 488.500 252.560 ;
 END
END B5
PIN B4
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER ME5 ;
  RECT 481.800 251.440 482.920 252.560 ;
  LAYER ME4 ;
  RECT 481.800 251.440 482.920 252.560 ;
  LAYER ME3 ;
  RECT 481.800 251.440 482.920 252.560 ;
  LAYER ME2 ;
  RECT 481.800 251.440 482.920 252.560 ;
  LAYER ME1 ;
  RECT 481.800 251.440 482.920 252.560 ;
 END
END B4
PIN B3
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER ME5 ;
  RECT 476.220 251.440 477.340 252.560 ;
  LAYER ME4 ;
  RECT 476.220 251.440 477.340 252.560 ;
  LAYER ME3 ;
  RECT 476.220 251.440 477.340 252.560 ;
  LAYER ME2 ;
  RECT 476.220 251.440 477.340 252.560 ;
  LAYER ME1 ;
  RECT 476.220 251.440 477.340 252.560 ;
 END
END B3
PIN B7
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER ME5 ;
  RECT 457.620 251.440 458.740 252.560 ;
  LAYER ME4 ;
  RECT 457.620 251.440 458.740 252.560 ;
  LAYER ME3 ;
  RECT 457.620 251.440 458.740 252.560 ;
  LAYER ME2 ;
  RECT 457.620 251.440 458.740 252.560 ;
  LAYER ME1 ;
  RECT 457.620 251.440 458.740 252.560 ;
 END
END B7
PIN B6
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER ME5 ;
  RECT 451.420 251.440 452.540 252.560 ;
  LAYER ME4 ;
  RECT 451.420 251.440 452.540 252.560 ;
  LAYER ME3 ;
  RECT 451.420 251.440 452.540 252.560 ;
  LAYER ME2 ;
  RECT 451.420 251.440 452.540 252.560 ;
  LAYER ME1 ;
  RECT 451.420 251.440 452.540 252.560 ;
 END
END B6
PIN DIB15
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER ME5 ;
  RECT 429.100 251.440 430.220 252.560 ;
  LAYER ME4 ;
  RECT 429.100 251.440 430.220 252.560 ;
  LAYER ME3 ;
  RECT 429.100 251.440 430.220 252.560 ;
  LAYER ME2 ;
  RECT 429.100 251.440 430.220 252.560 ;
  LAYER ME1 ;
  RECT 429.100 251.440 430.220 252.560 ;
 END
END DIB15
PIN DOB15
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME5 ;
  RECT 416.080 251.440 417.200 252.560 ;
  LAYER ME4 ;
  RECT 416.080 251.440 417.200 252.560 ;
  LAYER ME3 ;
  RECT 416.080 251.440 417.200 252.560 ;
  LAYER ME2 ;
  RECT 416.080 251.440 417.200 252.560 ;
  LAYER ME1 ;
  RECT 416.080 251.440 417.200 252.560 ;
 END
END DOB15
PIN DIB14
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER ME5 ;
  RECT 402.440 251.440 403.560 252.560 ;
  LAYER ME4 ;
  RECT 402.440 251.440 403.560 252.560 ;
  LAYER ME3 ;
  RECT 402.440 251.440 403.560 252.560 ;
  LAYER ME2 ;
  RECT 402.440 251.440 403.560 252.560 ;
  LAYER ME1 ;
  RECT 402.440 251.440 403.560 252.560 ;
 END
END DIB14
PIN DOB14
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME5 ;
  RECT 388.800 251.440 389.920 252.560 ;
  LAYER ME4 ;
  RECT 388.800 251.440 389.920 252.560 ;
  LAYER ME3 ;
  RECT 388.800 251.440 389.920 252.560 ;
  LAYER ME2 ;
  RECT 388.800 251.440 389.920 252.560 ;
  LAYER ME1 ;
  RECT 388.800 251.440 389.920 252.560 ;
 END
END DOB14
PIN DIB13
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER ME5 ;
  RECT 375.780 251.440 376.900 252.560 ;
  LAYER ME4 ;
  RECT 375.780 251.440 376.900 252.560 ;
  LAYER ME3 ;
  RECT 375.780 251.440 376.900 252.560 ;
  LAYER ME2 ;
  RECT 375.780 251.440 376.900 252.560 ;
  LAYER ME1 ;
  RECT 375.780 251.440 376.900 252.560 ;
 END
END DIB13
PIN DOB13
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME5 ;
  RECT 362.140 251.440 363.260 252.560 ;
  LAYER ME4 ;
  RECT 362.140 251.440 363.260 252.560 ;
  LAYER ME3 ;
  RECT 362.140 251.440 363.260 252.560 ;
  LAYER ME2 ;
  RECT 362.140 251.440 363.260 252.560 ;
  LAYER ME1 ;
  RECT 362.140 251.440 363.260 252.560 ;
 END
END DOB13
PIN DIB12
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER ME5 ;
  RECT 348.500 251.440 349.620 252.560 ;
  LAYER ME4 ;
  RECT 348.500 251.440 349.620 252.560 ;
  LAYER ME3 ;
  RECT 348.500 251.440 349.620 252.560 ;
  LAYER ME2 ;
  RECT 348.500 251.440 349.620 252.560 ;
  LAYER ME1 ;
  RECT 348.500 251.440 349.620 252.560 ;
 END
END DIB12
PIN DOB12
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME5 ;
  RECT 335.480 251.440 336.600 252.560 ;
  LAYER ME4 ;
  RECT 335.480 251.440 336.600 252.560 ;
  LAYER ME3 ;
  RECT 335.480 251.440 336.600 252.560 ;
  LAYER ME2 ;
  RECT 335.480 251.440 336.600 252.560 ;
  LAYER ME1 ;
  RECT 335.480 251.440 336.600 252.560 ;
 END
END DOB12
PIN DIB11
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER ME5 ;
  RECT 321.840 251.440 322.960 252.560 ;
  LAYER ME4 ;
  RECT 321.840 251.440 322.960 252.560 ;
  LAYER ME3 ;
  RECT 321.840 251.440 322.960 252.560 ;
  LAYER ME2 ;
  RECT 321.840 251.440 322.960 252.560 ;
  LAYER ME1 ;
  RECT 321.840 251.440 322.960 252.560 ;
 END
END DIB11
PIN DOB11
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME5 ;
  RECT 308.200 251.440 309.320 252.560 ;
  LAYER ME4 ;
  RECT 308.200 251.440 309.320 252.560 ;
  LAYER ME3 ;
  RECT 308.200 251.440 309.320 252.560 ;
  LAYER ME2 ;
  RECT 308.200 251.440 309.320 252.560 ;
  LAYER ME1 ;
  RECT 308.200 251.440 309.320 252.560 ;
 END
END DOB11
PIN DIB10
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER ME5 ;
  RECT 295.180 251.440 296.300 252.560 ;
  LAYER ME4 ;
  RECT 295.180 251.440 296.300 252.560 ;
  LAYER ME3 ;
  RECT 295.180 251.440 296.300 252.560 ;
  LAYER ME2 ;
  RECT 295.180 251.440 296.300 252.560 ;
  LAYER ME1 ;
  RECT 295.180 251.440 296.300 252.560 ;
 END
END DIB10
PIN DOB10
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME5 ;
  RECT 281.540 251.440 282.660 252.560 ;
  LAYER ME4 ;
  RECT 281.540 251.440 282.660 252.560 ;
  LAYER ME3 ;
  RECT 281.540 251.440 282.660 252.560 ;
  LAYER ME2 ;
  RECT 281.540 251.440 282.660 252.560 ;
  LAYER ME1 ;
  RECT 281.540 251.440 282.660 252.560 ;
 END
END DOB10
PIN DIB9
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER ME5 ;
  RECT 267.900 251.440 269.020 252.560 ;
  LAYER ME4 ;
  RECT 267.900 251.440 269.020 252.560 ;
  LAYER ME3 ;
  RECT 267.900 251.440 269.020 252.560 ;
  LAYER ME2 ;
  RECT 267.900 251.440 269.020 252.560 ;
  LAYER ME1 ;
  RECT 267.900 251.440 269.020 252.560 ;
 END
END DIB9
PIN DOB9
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME5 ;
  RECT 254.880 251.440 256.000 252.560 ;
  LAYER ME4 ;
  RECT 254.880 251.440 256.000 252.560 ;
  LAYER ME3 ;
  RECT 254.880 251.440 256.000 252.560 ;
  LAYER ME2 ;
  RECT 254.880 251.440 256.000 252.560 ;
  LAYER ME1 ;
  RECT 254.880 251.440 256.000 252.560 ;
 END
END DOB9
PIN DIB8
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER ME5 ;
  RECT 241.240 251.440 242.360 252.560 ;
  LAYER ME4 ;
  RECT 241.240 251.440 242.360 252.560 ;
  LAYER ME3 ;
  RECT 241.240 251.440 242.360 252.560 ;
  LAYER ME2 ;
  RECT 241.240 251.440 242.360 252.560 ;
  LAYER ME1 ;
  RECT 241.240 251.440 242.360 252.560 ;
 END
END DIB8
PIN DOB8
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME5 ;
  RECT 227.600 251.440 228.720 252.560 ;
  LAYER ME4 ;
  RECT 227.600 251.440 228.720 252.560 ;
  LAYER ME3 ;
  RECT 227.600 251.440 228.720 252.560 ;
  LAYER ME2 ;
  RECT 227.600 251.440 228.720 252.560 ;
  LAYER ME1 ;
  RECT 227.600 251.440 228.720 252.560 ;
 END
END DOB8
PIN DIB7
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER ME5 ;
  RECT 214.580 251.440 215.700 252.560 ;
  LAYER ME4 ;
  RECT 214.580 251.440 215.700 252.560 ;
  LAYER ME3 ;
  RECT 214.580 251.440 215.700 252.560 ;
  LAYER ME2 ;
  RECT 214.580 251.440 215.700 252.560 ;
  LAYER ME1 ;
  RECT 214.580 251.440 215.700 252.560 ;
 END
END DIB7
PIN DOB7
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME5 ;
  RECT 200.940 251.440 202.060 252.560 ;
  LAYER ME4 ;
  RECT 200.940 251.440 202.060 252.560 ;
  LAYER ME3 ;
  RECT 200.940 251.440 202.060 252.560 ;
  LAYER ME2 ;
  RECT 200.940 251.440 202.060 252.560 ;
  LAYER ME1 ;
  RECT 200.940 251.440 202.060 252.560 ;
 END
END DOB7
PIN DIB6
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER ME5 ;
  RECT 187.300 251.440 188.420 252.560 ;
  LAYER ME4 ;
  RECT 187.300 251.440 188.420 252.560 ;
  LAYER ME3 ;
  RECT 187.300 251.440 188.420 252.560 ;
  LAYER ME2 ;
  RECT 187.300 251.440 188.420 252.560 ;
  LAYER ME1 ;
  RECT 187.300 251.440 188.420 252.560 ;
 END
END DIB6
PIN DOB6
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME5 ;
  RECT 174.280 251.440 175.400 252.560 ;
  LAYER ME4 ;
  RECT 174.280 251.440 175.400 252.560 ;
  LAYER ME3 ;
  RECT 174.280 251.440 175.400 252.560 ;
  LAYER ME2 ;
  RECT 174.280 251.440 175.400 252.560 ;
  LAYER ME1 ;
  RECT 174.280 251.440 175.400 252.560 ;
 END
END DOB6
PIN DIB5
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER ME5 ;
  RECT 160.640 251.440 161.760 252.560 ;
  LAYER ME4 ;
  RECT 160.640 251.440 161.760 252.560 ;
  LAYER ME3 ;
  RECT 160.640 251.440 161.760 252.560 ;
  LAYER ME2 ;
  RECT 160.640 251.440 161.760 252.560 ;
  LAYER ME1 ;
  RECT 160.640 251.440 161.760 252.560 ;
 END
END DIB5
PIN DOB5
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME5 ;
  RECT 147.000 251.440 148.120 252.560 ;
  LAYER ME4 ;
  RECT 147.000 251.440 148.120 252.560 ;
  LAYER ME3 ;
  RECT 147.000 251.440 148.120 252.560 ;
  LAYER ME2 ;
  RECT 147.000 251.440 148.120 252.560 ;
  LAYER ME1 ;
  RECT 147.000 251.440 148.120 252.560 ;
 END
END DOB5
PIN DIB4
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER ME5 ;
  RECT 133.980 251.440 135.100 252.560 ;
  LAYER ME4 ;
  RECT 133.980 251.440 135.100 252.560 ;
  LAYER ME3 ;
  RECT 133.980 251.440 135.100 252.560 ;
  LAYER ME2 ;
  RECT 133.980 251.440 135.100 252.560 ;
  LAYER ME1 ;
  RECT 133.980 251.440 135.100 252.560 ;
 END
END DIB4
PIN DOB4
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME5 ;
  RECT 120.340 251.440 121.460 252.560 ;
  LAYER ME4 ;
  RECT 120.340 251.440 121.460 252.560 ;
  LAYER ME3 ;
  RECT 120.340 251.440 121.460 252.560 ;
  LAYER ME2 ;
  RECT 120.340 251.440 121.460 252.560 ;
  LAYER ME1 ;
  RECT 120.340 251.440 121.460 252.560 ;
 END
END DOB4
PIN DIB3
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER ME5 ;
  RECT 106.700 251.440 107.820 252.560 ;
  LAYER ME4 ;
  RECT 106.700 251.440 107.820 252.560 ;
  LAYER ME3 ;
  RECT 106.700 251.440 107.820 252.560 ;
  LAYER ME2 ;
  RECT 106.700 251.440 107.820 252.560 ;
  LAYER ME1 ;
  RECT 106.700 251.440 107.820 252.560 ;
 END
END DIB3
PIN DOB3
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME5 ;
  RECT 93.680 251.440 94.800 252.560 ;
  LAYER ME4 ;
  RECT 93.680 251.440 94.800 252.560 ;
  LAYER ME3 ;
  RECT 93.680 251.440 94.800 252.560 ;
  LAYER ME2 ;
  RECT 93.680 251.440 94.800 252.560 ;
  LAYER ME1 ;
  RECT 93.680 251.440 94.800 252.560 ;
 END
END DOB3
PIN DIB2
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER ME5 ;
  RECT 80.040 251.440 81.160 252.560 ;
  LAYER ME4 ;
  RECT 80.040 251.440 81.160 252.560 ;
  LAYER ME3 ;
  RECT 80.040 251.440 81.160 252.560 ;
  LAYER ME2 ;
  RECT 80.040 251.440 81.160 252.560 ;
  LAYER ME1 ;
  RECT 80.040 251.440 81.160 252.560 ;
 END
END DIB2
PIN DOB2
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME5 ;
  RECT 66.400 251.440 67.520 252.560 ;
  LAYER ME4 ;
  RECT 66.400 251.440 67.520 252.560 ;
  LAYER ME3 ;
  RECT 66.400 251.440 67.520 252.560 ;
  LAYER ME2 ;
  RECT 66.400 251.440 67.520 252.560 ;
  LAYER ME1 ;
  RECT 66.400 251.440 67.520 252.560 ;
 END
END DOB2
PIN DIB1
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER ME5 ;
  RECT 52.760 251.440 53.880 252.560 ;
  LAYER ME4 ;
  RECT 52.760 251.440 53.880 252.560 ;
  LAYER ME3 ;
  RECT 52.760 251.440 53.880 252.560 ;
  LAYER ME2 ;
  RECT 52.760 251.440 53.880 252.560 ;
  LAYER ME1 ;
  RECT 52.760 251.440 53.880 252.560 ;
 END
END DIB1
PIN DOB1
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME5 ;
  RECT 39.740 251.440 40.860 252.560 ;
  LAYER ME4 ;
  RECT 39.740 251.440 40.860 252.560 ;
  LAYER ME3 ;
  RECT 39.740 251.440 40.860 252.560 ;
  LAYER ME2 ;
  RECT 39.740 251.440 40.860 252.560 ;
  LAYER ME1 ;
  RECT 39.740 251.440 40.860 252.560 ;
 END
END DOB1
PIN DIB0
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER ME5 ;
  RECT 26.100 251.440 27.220 252.560 ;
  LAYER ME4 ;
  RECT 26.100 251.440 27.220 252.560 ;
  LAYER ME3 ;
  RECT 26.100 251.440 27.220 252.560 ;
  LAYER ME2 ;
  RECT 26.100 251.440 27.220 252.560 ;
  LAYER ME1 ;
  RECT 26.100 251.440 27.220 252.560 ;
 END
END DIB0
PIN DOB0
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME5 ;
  RECT 12.460 251.440 13.580 252.560 ;
  LAYER ME4 ;
  RECT 12.460 251.440 13.580 252.560 ;
  LAYER ME3 ;
  RECT 12.460 251.440 13.580 252.560 ;
  LAYER ME2 ;
  RECT 12.460 251.440 13.580 252.560 ;
  LAYER ME1 ;
  RECT 12.460 251.440 13.580 252.560 ;
 END
END DOB0
PIN DIA31
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER ME5 ;
  RECT 949.900 0.000 951.020 1.120 ;
  LAYER ME4 ;
  RECT 949.900 0.000 951.020 1.120 ;
  LAYER ME3 ;
  RECT 949.900 0.000 951.020 1.120 ;
  LAYER ME2 ;
  RECT 949.900 0.000 951.020 1.120 ;
  LAYER ME1 ;
  RECT 949.900 0.000 951.020 1.120 ;
 END
END DIA31
PIN DOA31
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER ME5 ;
  RECT 936.260 0.000 937.380 1.120 ;
  LAYER ME4 ;
  RECT 936.260 0.000 937.380 1.120 ;
  LAYER ME3 ;
  RECT 936.260 0.000 937.380 1.120 ;
  LAYER ME2 ;
  RECT 936.260 0.000 937.380 1.120 ;
  LAYER ME1 ;
  RECT 936.260 0.000 937.380 1.120 ;
 END
END DOA31
PIN DIA30
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER ME5 ;
  RECT 923.240 0.000 924.360 1.120 ;
  LAYER ME4 ;
  RECT 923.240 0.000 924.360 1.120 ;
  LAYER ME3 ;
  RECT 923.240 0.000 924.360 1.120 ;
  LAYER ME2 ;
  RECT 923.240 0.000 924.360 1.120 ;
  LAYER ME1 ;
  RECT 923.240 0.000 924.360 1.120 ;
 END
END DIA30
PIN DOA30
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME5 ;
  RECT 909.600 0.000 910.720 1.120 ;
  LAYER ME4 ;
  RECT 909.600 0.000 910.720 1.120 ;
  LAYER ME3 ;
  RECT 909.600 0.000 910.720 1.120 ;
  LAYER ME2 ;
  RECT 909.600 0.000 910.720 1.120 ;
  LAYER ME1 ;
  RECT 909.600 0.000 910.720 1.120 ;
 END
END DOA30
PIN DIA29
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER ME5 ;
  RECT 895.960 0.000 897.080 1.120 ;
  LAYER ME4 ;
  RECT 895.960 0.000 897.080 1.120 ;
  LAYER ME3 ;
  RECT 895.960 0.000 897.080 1.120 ;
  LAYER ME2 ;
  RECT 895.960 0.000 897.080 1.120 ;
  LAYER ME1 ;
  RECT 895.960 0.000 897.080 1.120 ;
 END
END DIA29
PIN DOA29
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER ME5 ;
  RECT 882.940 0.000 884.060 1.120 ;
  LAYER ME4 ;
  RECT 882.940 0.000 884.060 1.120 ;
  LAYER ME3 ;
  RECT 882.940 0.000 884.060 1.120 ;
  LAYER ME2 ;
  RECT 882.940 0.000 884.060 1.120 ;
  LAYER ME1 ;
  RECT 882.940 0.000 884.060 1.120 ;
 END
END DOA29
PIN DIA28
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER ME5 ;
  RECT 869.300 0.000 870.420 1.120 ;
  LAYER ME4 ;
  RECT 869.300 0.000 870.420 1.120 ;
  LAYER ME3 ;
  RECT 869.300 0.000 870.420 1.120 ;
  LAYER ME2 ;
  RECT 869.300 0.000 870.420 1.120 ;
  LAYER ME1 ;
  RECT 869.300 0.000 870.420 1.120 ;
 END
END DIA28
PIN DOA28
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME5 ;
  RECT 855.660 0.000 856.780 1.120 ;
  LAYER ME4 ;
  RECT 855.660 0.000 856.780 1.120 ;
  LAYER ME3 ;
  RECT 855.660 0.000 856.780 1.120 ;
  LAYER ME2 ;
  RECT 855.660 0.000 856.780 1.120 ;
  LAYER ME1 ;
  RECT 855.660 0.000 856.780 1.120 ;
 END
END DOA28
PIN DIA27
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER ME5 ;
  RECT 842.640 0.000 843.760 1.120 ;
  LAYER ME4 ;
  RECT 842.640 0.000 843.760 1.120 ;
  LAYER ME3 ;
  RECT 842.640 0.000 843.760 1.120 ;
  LAYER ME2 ;
  RECT 842.640 0.000 843.760 1.120 ;
  LAYER ME1 ;
  RECT 842.640 0.000 843.760 1.120 ;
 END
END DIA27
PIN DOA27
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME5 ;
  RECT 829.000 0.000 830.120 1.120 ;
  LAYER ME4 ;
  RECT 829.000 0.000 830.120 1.120 ;
  LAYER ME3 ;
  RECT 829.000 0.000 830.120 1.120 ;
  LAYER ME2 ;
  RECT 829.000 0.000 830.120 1.120 ;
  LAYER ME1 ;
  RECT 829.000 0.000 830.120 1.120 ;
 END
END DOA27
PIN DIA26
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER ME5 ;
  RECT 815.360 0.000 816.480 1.120 ;
  LAYER ME4 ;
  RECT 815.360 0.000 816.480 1.120 ;
  LAYER ME3 ;
  RECT 815.360 0.000 816.480 1.120 ;
  LAYER ME2 ;
  RECT 815.360 0.000 816.480 1.120 ;
  LAYER ME1 ;
  RECT 815.360 0.000 816.480 1.120 ;
 END
END DIA26
PIN DOA26
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER ME5 ;
  RECT 802.340 0.000 803.460 1.120 ;
  LAYER ME4 ;
  RECT 802.340 0.000 803.460 1.120 ;
  LAYER ME3 ;
  RECT 802.340 0.000 803.460 1.120 ;
  LAYER ME2 ;
  RECT 802.340 0.000 803.460 1.120 ;
  LAYER ME1 ;
  RECT 802.340 0.000 803.460 1.120 ;
 END
END DOA26
PIN DIA25
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER ME5 ;
  RECT 788.700 0.000 789.820 1.120 ;
  LAYER ME4 ;
  RECT 788.700 0.000 789.820 1.120 ;
  LAYER ME3 ;
  RECT 788.700 0.000 789.820 1.120 ;
  LAYER ME2 ;
  RECT 788.700 0.000 789.820 1.120 ;
  LAYER ME1 ;
  RECT 788.700 0.000 789.820 1.120 ;
 END
END DIA25
PIN DOA25
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME5 ;
  RECT 775.060 0.000 776.180 1.120 ;
  LAYER ME4 ;
  RECT 775.060 0.000 776.180 1.120 ;
  LAYER ME3 ;
  RECT 775.060 0.000 776.180 1.120 ;
  LAYER ME2 ;
  RECT 775.060 0.000 776.180 1.120 ;
  LAYER ME1 ;
  RECT 775.060 0.000 776.180 1.120 ;
 END
END DOA25
PIN DIA24
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER ME5 ;
  RECT 761.420 0.000 762.540 1.120 ;
  LAYER ME4 ;
  RECT 761.420 0.000 762.540 1.120 ;
  LAYER ME3 ;
  RECT 761.420 0.000 762.540 1.120 ;
  LAYER ME2 ;
  RECT 761.420 0.000 762.540 1.120 ;
  LAYER ME1 ;
  RECT 761.420 0.000 762.540 1.120 ;
 END
END DIA24
PIN DOA24
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME5 ;
  RECT 748.400 0.000 749.520 1.120 ;
  LAYER ME4 ;
  RECT 748.400 0.000 749.520 1.120 ;
  LAYER ME3 ;
  RECT 748.400 0.000 749.520 1.120 ;
  LAYER ME2 ;
  RECT 748.400 0.000 749.520 1.120 ;
  LAYER ME1 ;
  RECT 748.400 0.000 749.520 1.120 ;
 END
END DOA24
PIN DIA23
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER ME5 ;
  RECT 734.760 0.000 735.880 1.120 ;
  LAYER ME4 ;
  RECT 734.760 0.000 735.880 1.120 ;
  LAYER ME3 ;
  RECT 734.760 0.000 735.880 1.120 ;
  LAYER ME2 ;
  RECT 734.760 0.000 735.880 1.120 ;
  LAYER ME1 ;
  RECT 734.760 0.000 735.880 1.120 ;
 END
END DIA23
PIN DOA23
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER ME5 ;
  RECT 721.120 0.000 722.240 1.120 ;
  LAYER ME4 ;
  RECT 721.120 0.000 722.240 1.120 ;
  LAYER ME3 ;
  RECT 721.120 0.000 722.240 1.120 ;
  LAYER ME2 ;
  RECT 721.120 0.000 722.240 1.120 ;
  LAYER ME1 ;
  RECT 721.120 0.000 722.240 1.120 ;
 END
END DOA23
PIN DIA22
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER ME5 ;
  RECT 708.100 0.000 709.220 1.120 ;
  LAYER ME4 ;
  RECT 708.100 0.000 709.220 1.120 ;
  LAYER ME3 ;
  RECT 708.100 0.000 709.220 1.120 ;
  LAYER ME2 ;
  RECT 708.100 0.000 709.220 1.120 ;
  LAYER ME1 ;
  RECT 708.100 0.000 709.220 1.120 ;
 END
END DIA22
PIN DOA22
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME5 ;
  RECT 694.460 0.000 695.580 1.120 ;
  LAYER ME4 ;
  RECT 694.460 0.000 695.580 1.120 ;
  LAYER ME3 ;
  RECT 694.460 0.000 695.580 1.120 ;
  LAYER ME2 ;
  RECT 694.460 0.000 695.580 1.120 ;
  LAYER ME1 ;
  RECT 694.460 0.000 695.580 1.120 ;
 END
END DOA22
PIN DIA21
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER ME5 ;
  RECT 680.820 0.000 681.940 1.120 ;
  LAYER ME4 ;
  RECT 680.820 0.000 681.940 1.120 ;
  LAYER ME3 ;
  RECT 680.820 0.000 681.940 1.120 ;
  LAYER ME2 ;
  RECT 680.820 0.000 681.940 1.120 ;
  LAYER ME1 ;
  RECT 680.820 0.000 681.940 1.120 ;
 END
END DIA21
PIN DOA21
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER ME5 ;
  RECT 667.800 0.000 668.920 1.120 ;
  LAYER ME4 ;
  RECT 667.800 0.000 668.920 1.120 ;
  LAYER ME3 ;
  RECT 667.800 0.000 668.920 1.120 ;
  LAYER ME2 ;
  RECT 667.800 0.000 668.920 1.120 ;
  LAYER ME1 ;
  RECT 667.800 0.000 668.920 1.120 ;
 END
END DOA21
PIN DIA20
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER ME5 ;
  RECT 654.160 0.000 655.280 1.120 ;
  LAYER ME4 ;
  RECT 654.160 0.000 655.280 1.120 ;
  LAYER ME3 ;
  RECT 654.160 0.000 655.280 1.120 ;
  LAYER ME2 ;
  RECT 654.160 0.000 655.280 1.120 ;
  LAYER ME1 ;
  RECT 654.160 0.000 655.280 1.120 ;
 END
END DIA20
PIN DOA20
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER ME5 ;
  RECT 640.520 0.000 641.640 1.120 ;
  LAYER ME4 ;
  RECT 640.520 0.000 641.640 1.120 ;
  LAYER ME3 ;
  RECT 640.520 0.000 641.640 1.120 ;
  LAYER ME2 ;
  RECT 640.520 0.000 641.640 1.120 ;
  LAYER ME1 ;
  RECT 640.520 0.000 641.640 1.120 ;
 END
END DOA20
PIN DIA19
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER ME5 ;
  RECT 627.500 0.000 628.620 1.120 ;
  LAYER ME4 ;
  RECT 627.500 0.000 628.620 1.120 ;
  LAYER ME3 ;
  RECT 627.500 0.000 628.620 1.120 ;
  LAYER ME2 ;
  RECT 627.500 0.000 628.620 1.120 ;
  LAYER ME1 ;
  RECT 627.500 0.000 628.620 1.120 ;
 END
END DIA19
PIN DOA19
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME5 ;
  RECT 613.860 0.000 614.980 1.120 ;
  LAYER ME4 ;
  RECT 613.860 0.000 614.980 1.120 ;
  LAYER ME3 ;
  RECT 613.860 0.000 614.980 1.120 ;
  LAYER ME2 ;
  RECT 613.860 0.000 614.980 1.120 ;
  LAYER ME1 ;
  RECT 613.860 0.000 614.980 1.120 ;
 END
END DOA19
PIN DIA18
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER ME5 ;
  RECT 600.220 0.000 601.340 1.120 ;
  LAYER ME4 ;
  RECT 600.220 0.000 601.340 1.120 ;
  LAYER ME3 ;
  RECT 600.220 0.000 601.340 1.120 ;
  LAYER ME2 ;
  RECT 600.220 0.000 601.340 1.120 ;
  LAYER ME1 ;
  RECT 600.220 0.000 601.340 1.120 ;
 END
END DIA18
PIN DOA18
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER ME5 ;
  RECT 587.200 0.000 588.320 1.120 ;
  LAYER ME4 ;
  RECT 587.200 0.000 588.320 1.120 ;
  LAYER ME3 ;
  RECT 587.200 0.000 588.320 1.120 ;
  LAYER ME2 ;
  RECT 587.200 0.000 588.320 1.120 ;
  LAYER ME1 ;
  RECT 587.200 0.000 588.320 1.120 ;
 END
END DOA18
PIN DIA17
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER ME5 ;
  RECT 573.560 0.000 574.680 1.120 ;
  LAYER ME4 ;
  RECT 573.560 0.000 574.680 1.120 ;
  LAYER ME3 ;
  RECT 573.560 0.000 574.680 1.120 ;
  LAYER ME2 ;
  RECT 573.560 0.000 574.680 1.120 ;
  LAYER ME1 ;
  RECT 573.560 0.000 574.680 1.120 ;
 END
END DIA17
PIN DOA17
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER ME5 ;
  RECT 559.920 0.000 561.040 1.120 ;
  LAYER ME4 ;
  RECT 559.920 0.000 561.040 1.120 ;
  LAYER ME3 ;
  RECT 559.920 0.000 561.040 1.120 ;
  LAYER ME2 ;
  RECT 559.920 0.000 561.040 1.120 ;
  LAYER ME1 ;
  RECT 559.920 0.000 561.040 1.120 ;
 END
END DOA17
PIN DIA16
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER ME5 ;
  RECT 546.900 0.000 548.020 1.120 ;
  LAYER ME4 ;
  RECT 546.900 0.000 548.020 1.120 ;
  LAYER ME3 ;
  RECT 546.900 0.000 548.020 1.120 ;
  LAYER ME2 ;
  RECT 546.900 0.000 548.020 1.120 ;
  LAYER ME1 ;
  RECT 546.900 0.000 548.020 1.120 ;
 END
END DIA16
PIN DOA16
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME5 ;
  RECT 533.260 0.000 534.380 1.120 ;
  LAYER ME4 ;
  RECT 533.260 0.000 534.380 1.120 ;
  LAYER ME3 ;
  RECT 533.260 0.000 534.380 1.120 ;
  LAYER ME2 ;
  RECT 533.260 0.000 534.380 1.120 ;
  LAYER ME1 ;
  RECT 533.260 0.000 534.380 1.120 ;
 END
END DOA16
PIN CKA
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER ME5 ;
  RECT 511.560 0.000 512.680 1.120 ;
  LAYER ME4 ;
  RECT 511.560 0.000 512.680 1.120 ;
  LAYER ME3 ;
  RECT 511.560 0.000 512.680 1.120 ;
  LAYER ME2 ;
  RECT 511.560 0.000 512.680 1.120 ;
  LAYER ME1 ;
  RECT 511.560 0.000 512.680 1.120 ;
 END
END CKA
PIN CSA
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER ME5 ;
  RECT 509.080 0.000 510.200 1.120 ;
  LAYER ME4 ;
  RECT 509.080 0.000 510.200 1.120 ;
  LAYER ME3 ;
  RECT 509.080 0.000 510.200 1.120 ;
  LAYER ME2 ;
  RECT 509.080 0.000 510.200 1.120 ;
  LAYER ME1 ;
  RECT 509.080 0.000 510.200 1.120 ;
 END
END CSA
PIN WEAN
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER ME5 ;
  RECT 507.220 0.000 508.340 1.120 ;
  LAYER ME4 ;
  RECT 507.220 0.000 508.340 1.120 ;
  LAYER ME3 ;
  RECT 507.220 0.000 508.340 1.120 ;
  LAYER ME2 ;
  RECT 507.220 0.000 508.340 1.120 ;
  LAYER ME1 ;
  RECT 507.220 0.000 508.340 1.120 ;
 END
END WEAN
PIN A2
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER ME5 ;
  RECT 503.500 0.000 504.620 1.120 ;
  LAYER ME4 ;
  RECT 503.500 0.000 504.620 1.120 ;
  LAYER ME3 ;
  RECT 503.500 0.000 504.620 1.120 ;
  LAYER ME2 ;
  RECT 503.500 0.000 504.620 1.120 ;
  LAYER ME1 ;
  RECT 503.500 0.000 504.620 1.120 ;
 END
END A2
PIN OEA
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER ME5 ;
  RECT 499.780 0.000 500.900 1.120 ;
  LAYER ME4 ;
  RECT 499.780 0.000 500.900 1.120 ;
  LAYER ME3 ;
  RECT 499.780 0.000 500.900 1.120 ;
  LAYER ME2 ;
  RECT 499.780 0.000 500.900 1.120 ;
  LAYER ME1 ;
  RECT 499.780 0.000 500.900 1.120 ;
 END
END OEA
PIN A1
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER ME5 ;
  RECT 497.920 0.000 499.040 1.120 ;
  LAYER ME4 ;
  RECT 497.920 0.000 499.040 1.120 ;
  LAYER ME3 ;
  RECT 497.920 0.000 499.040 1.120 ;
  LAYER ME2 ;
  RECT 497.920 0.000 499.040 1.120 ;
  LAYER ME1 ;
  RECT 497.920 0.000 499.040 1.120 ;
 END
END A1
PIN A0
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER ME5 ;
  RECT 496.060 0.000 497.180 1.120 ;
  LAYER ME4 ;
  RECT 496.060 0.000 497.180 1.120 ;
  LAYER ME3 ;
  RECT 496.060 0.000 497.180 1.120 ;
  LAYER ME2 ;
  RECT 496.060 0.000 497.180 1.120 ;
  LAYER ME1 ;
  RECT 496.060 0.000 497.180 1.120 ;
 END
END A0
PIN A5
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER ME5 ;
  RECT 487.380 0.000 488.500 1.120 ;
  LAYER ME4 ;
  RECT 487.380 0.000 488.500 1.120 ;
  LAYER ME3 ;
  RECT 487.380 0.000 488.500 1.120 ;
  LAYER ME2 ;
  RECT 487.380 0.000 488.500 1.120 ;
  LAYER ME1 ;
  RECT 487.380 0.000 488.500 1.120 ;
 END
END A5
PIN A4
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER ME5 ;
  RECT 481.800 0.000 482.920 1.120 ;
  LAYER ME4 ;
  RECT 481.800 0.000 482.920 1.120 ;
  LAYER ME3 ;
  RECT 481.800 0.000 482.920 1.120 ;
  LAYER ME2 ;
  RECT 481.800 0.000 482.920 1.120 ;
  LAYER ME1 ;
  RECT 481.800 0.000 482.920 1.120 ;
 END
END A4
PIN A3
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER ME5 ;
  RECT 476.220 0.000 477.340 1.120 ;
  LAYER ME4 ;
  RECT 476.220 0.000 477.340 1.120 ;
  LAYER ME3 ;
  RECT 476.220 0.000 477.340 1.120 ;
  LAYER ME2 ;
  RECT 476.220 0.000 477.340 1.120 ;
  LAYER ME1 ;
  RECT 476.220 0.000 477.340 1.120 ;
 END
END A3
PIN A7
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER ME5 ;
  RECT 457.620 0.000 458.740 1.120 ;
  LAYER ME4 ;
  RECT 457.620 0.000 458.740 1.120 ;
  LAYER ME3 ;
  RECT 457.620 0.000 458.740 1.120 ;
  LAYER ME2 ;
  RECT 457.620 0.000 458.740 1.120 ;
  LAYER ME1 ;
  RECT 457.620 0.000 458.740 1.120 ;
 END
END A7
PIN A6
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER ME5 ;
  RECT 451.420 0.000 452.540 1.120 ;
  LAYER ME4 ;
  RECT 451.420 0.000 452.540 1.120 ;
  LAYER ME3 ;
  RECT 451.420 0.000 452.540 1.120 ;
  LAYER ME2 ;
  RECT 451.420 0.000 452.540 1.120 ;
  LAYER ME1 ;
  RECT 451.420 0.000 452.540 1.120 ;
 END
END A6
PIN DIA15
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER ME5 ;
  RECT 429.100 0.000 430.220 1.120 ;
  LAYER ME4 ;
  RECT 429.100 0.000 430.220 1.120 ;
  LAYER ME3 ;
  RECT 429.100 0.000 430.220 1.120 ;
  LAYER ME2 ;
  RECT 429.100 0.000 430.220 1.120 ;
  LAYER ME1 ;
  RECT 429.100 0.000 430.220 1.120 ;
 END
END DIA15
PIN DOA15
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME5 ;
  RECT 416.080 0.000 417.200 1.120 ;
  LAYER ME4 ;
  RECT 416.080 0.000 417.200 1.120 ;
  LAYER ME3 ;
  RECT 416.080 0.000 417.200 1.120 ;
  LAYER ME2 ;
  RECT 416.080 0.000 417.200 1.120 ;
  LAYER ME1 ;
  RECT 416.080 0.000 417.200 1.120 ;
 END
END DOA15
PIN DIA14
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER ME5 ;
  RECT 402.440 0.000 403.560 1.120 ;
  LAYER ME4 ;
  RECT 402.440 0.000 403.560 1.120 ;
  LAYER ME3 ;
  RECT 402.440 0.000 403.560 1.120 ;
  LAYER ME2 ;
  RECT 402.440 0.000 403.560 1.120 ;
  LAYER ME1 ;
  RECT 402.440 0.000 403.560 1.120 ;
 END
END DIA14
PIN DOA14
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER ME5 ;
  RECT 388.800 0.000 389.920 1.120 ;
  LAYER ME4 ;
  RECT 388.800 0.000 389.920 1.120 ;
  LAYER ME3 ;
  RECT 388.800 0.000 389.920 1.120 ;
  LAYER ME2 ;
  RECT 388.800 0.000 389.920 1.120 ;
  LAYER ME1 ;
  RECT 388.800 0.000 389.920 1.120 ;
 END
END DOA14
PIN DIA13
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER ME5 ;
  RECT 375.780 0.000 376.900 1.120 ;
  LAYER ME4 ;
  RECT 375.780 0.000 376.900 1.120 ;
  LAYER ME3 ;
  RECT 375.780 0.000 376.900 1.120 ;
  LAYER ME2 ;
  RECT 375.780 0.000 376.900 1.120 ;
  LAYER ME1 ;
  RECT 375.780 0.000 376.900 1.120 ;
 END
END DIA13
PIN DOA13
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME5 ;
  RECT 362.140 0.000 363.260 1.120 ;
  LAYER ME4 ;
  RECT 362.140 0.000 363.260 1.120 ;
  LAYER ME3 ;
  RECT 362.140 0.000 363.260 1.120 ;
  LAYER ME2 ;
  RECT 362.140 0.000 363.260 1.120 ;
  LAYER ME1 ;
  RECT 362.140 0.000 363.260 1.120 ;
 END
END DOA13
PIN DIA12
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER ME5 ;
  RECT 348.500 0.000 349.620 1.120 ;
  LAYER ME4 ;
  RECT 348.500 0.000 349.620 1.120 ;
  LAYER ME3 ;
  RECT 348.500 0.000 349.620 1.120 ;
  LAYER ME2 ;
  RECT 348.500 0.000 349.620 1.120 ;
  LAYER ME1 ;
  RECT 348.500 0.000 349.620 1.120 ;
 END
END DIA12
PIN DOA12
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER ME5 ;
  RECT 335.480 0.000 336.600 1.120 ;
  LAYER ME4 ;
  RECT 335.480 0.000 336.600 1.120 ;
  LAYER ME3 ;
  RECT 335.480 0.000 336.600 1.120 ;
  LAYER ME2 ;
  RECT 335.480 0.000 336.600 1.120 ;
  LAYER ME1 ;
  RECT 335.480 0.000 336.600 1.120 ;
 END
END DOA12
PIN DIA11
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER ME5 ;
  RECT 321.840 0.000 322.960 1.120 ;
  LAYER ME4 ;
  RECT 321.840 0.000 322.960 1.120 ;
  LAYER ME3 ;
  RECT 321.840 0.000 322.960 1.120 ;
  LAYER ME2 ;
  RECT 321.840 0.000 322.960 1.120 ;
  LAYER ME1 ;
  RECT 321.840 0.000 322.960 1.120 ;
 END
END DIA11
PIN DOA11
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER ME5 ;
  RECT 308.200 0.000 309.320 1.120 ;
  LAYER ME4 ;
  RECT 308.200 0.000 309.320 1.120 ;
  LAYER ME3 ;
  RECT 308.200 0.000 309.320 1.120 ;
  LAYER ME2 ;
  RECT 308.200 0.000 309.320 1.120 ;
  LAYER ME1 ;
  RECT 308.200 0.000 309.320 1.120 ;
 END
END DOA11
PIN DIA10
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER ME5 ;
  RECT 295.180 0.000 296.300 1.120 ;
  LAYER ME4 ;
  RECT 295.180 0.000 296.300 1.120 ;
  LAYER ME3 ;
  RECT 295.180 0.000 296.300 1.120 ;
  LAYER ME2 ;
  RECT 295.180 0.000 296.300 1.120 ;
  LAYER ME1 ;
  RECT 295.180 0.000 296.300 1.120 ;
 END
END DIA10
PIN DOA10
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME5 ;
  RECT 281.540 0.000 282.660 1.120 ;
  LAYER ME4 ;
  RECT 281.540 0.000 282.660 1.120 ;
  LAYER ME3 ;
  RECT 281.540 0.000 282.660 1.120 ;
  LAYER ME2 ;
  RECT 281.540 0.000 282.660 1.120 ;
  LAYER ME1 ;
  RECT 281.540 0.000 282.660 1.120 ;
 END
END DOA10
PIN DIA9
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER ME5 ;
  RECT 267.900 0.000 269.020 1.120 ;
  LAYER ME4 ;
  RECT 267.900 0.000 269.020 1.120 ;
  LAYER ME3 ;
  RECT 267.900 0.000 269.020 1.120 ;
  LAYER ME2 ;
  RECT 267.900 0.000 269.020 1.120 ;
  LAYER ME1 ;
  RECT 267.900 0.000 269.020 1.120 ;
 END
END DIA9
PIN DOA9
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER ME5 ;
  RECT 254.880 0.000 256.000 1.120 ;
  LAYER ME4 ;
  RECT 254.880 0.000 256.000 1.120 ;
  LAYER ME3 ;
  RECT 254.880 0.000 256.000 1.120 ;
  LAYER ME2 ;
  RECT 254.880 0.000 256.000 1.120 ;
  LAYER ME1 ;
  RECT 254.880 0.000 256.000 1.120 ;
 END
END DOA9
PIN DIA8
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER ME5 ;
  RECT 241.240 0.000 242.360 1.120 ;
  LAYER ME4 ;
  RECT 241.240 0.000 242.360 1.120 ;
  LAYER ME3 ;
  RECT 241.240 0.000 242.360 1.120 ;
  LAYER ME2 ;
  RECT 241.240 0.000 242.360 1.120 ;
  LAYER ME1 ;
  RECT 241.240 0.000 242.360 1.120 ;
 END
END DIA8
PIN DOA8
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER ME5 ;
  RECT 227.600 0.000 228.720 1.120 ;
  LAYER ME4 ;
  RECT 227.600 0.000 228.720 1.120 ;
  LAYER ME3 ;
  RECT 227.600 0.000 228.720 1.120 ;
  LAYER ME2 ;
  RECT 227.600 0.000 228.720 1.120 ;
  LAYER ME1 ;
  RECT 227.600 0.000 228.720 1.120 ;
 END
END DOA8
PIN DIA7
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER ME5 ;
  RECT 214.580 0.000 215.700 1.120 ;
  LAYER ME4 ;
  RECT 214.580 0.000 215.700 1.120 ;
  LAYER ME3 ;
  RECT 214.580 0.000 215.700 1.120 ;
  LAYER ME2 ;
  RECT 214.580 0.000 215.700 1.120 ;
  LAYER ME1 ;
  RECT 214.580 0.000 215.700 1.120 ;
 END
END DIA7
PIN DOA7
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME5 ;
  RECT 200.940 0.000 202.060 1.120 ;
  LAYER ME4 ;
  RECT 200.940 0.000 202.060 1.120 ;
  LAYER ME3 ;
  RECT 200.940 0.000 202.060 1.120 ;
  LAYER ME2 ;
  RECT 200.940 0.000 202.060 1.120 ;
  LAYER ME1 ;
  RECT 200.940 0.000 202.060 1.120 ;
 END
END DOA7
PIN DIA6
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER ME5 ;
  RECT 187.300 0.000 188.420 1.120 ;
  LAYER ME4 ;
  RECT 187.300 0.000 188.420 1.120 ;
  LAYER ME3 ;
  RECT 187.300 0.000 188.420 1.120 ;
  LAYER ME2 ;
  RECT 187.300 0.000 188.420 1.120 ;
  LAYER ME1 ;
  RECT 187.300 0.000 188.420 1.120 ;
 END
END DIA6
PIN DOA6
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER ME5 ;
  RECT 174.280 0.000 175.400 1.120 ;
  LAYER ME4 ;
  RECT 174.280 0.000 175.400 1.120 ;
  LAYER ME3 ;
  RECT 174.280 0.000 175.400 1.120 ;
  LAYER ME2 ;
  RECT 174.280 0.000 175.400 1.120 ;
  LAYER ME1 ;
  RECT 174.280 0.000 175.400 1.120 ;
 END
END DOA6
PIN DIA5
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER ME5 ;
  RECT 160.640 0.000 161.760 1.120 ;
  LAYER ME4 ;
  RECT 160.640 0.000 161.760 1.120 ;
  LAYER ME3 ;
  RECT 160.640 0.000 161.760 1.120 ;
  LAYER ME2 ;
  RECT 160.640 0.000 161.760 1.120 ;
  LAYER ME1 ;
  RECT 160.640 0.000 161.760 1.120 ;
 END
END DIA5
PIN DOA5
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER ME5 ;
  RECT 147.000 0.000 148.120 1.120 ;
  LAYER ME4 ;
  RECT 147.000 0.000 148.120 1.120 ;
  LAYER ME3 ;
  RECT 147.000 0.000 148.120 1.120 ;
  LAYER ME2 ;
  RECT 147.000 0.000 148.120 1.120 ;
  LAYER ME1 ;
  RECT 147.000 0.000 148.120 1.120 ;
 END
END DOA5
PIN DIA4
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER ME5 ;
  RECT 133.980 0.000 135.100 1.120 ;
  LAYER ME4 ;
  RECT 133.980 0.000 135.100 1.120 ;
  LAYER ME3 ;
  RECT 133.980 0.000 135.100 1.120 ;
  LAYER ME2 ;
  RECT 133.980 0.000 135.100 1.120 ;
  LAYER ME1 ;
  RECT 133.980 0.000 135.100 1.120 ;
 END
END DIA4
PIN DOA4
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME5 ;
  RECT 120.340 0.000 121.460 1.120 ;
  LAYER ME4 ;
  RECT 120.340 0.000 121.460 1.120 ;
  LAYER ME3 ;
  RECT 120.340 0.000 121.460 1.120 ;
  LAYER ME2 ;
  RECT 120.340 0.000 121.460 1.120 ;
  LAYER ME1 ;
  RECT 120.340 0.000 121.460 1.120 ;
 END
END DOA4
PIN DIA3
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER ME5 ;
  RECT 106.700 0.000 107.820 1.120 ;
  LAYER ME4 ;
  RECT 106.700 0.000 107.820 1.120 ;
  LAYER ME3 ;
  RECT 106.700 0.000 107.820 1.120 ;
  LAYER ME2 ;
  RECT 106.700 0.000 107.820 1.120 ;
  LAYER ME1 ;
  RECT 106.700 0.000 107.820 1.120 ;
 END
END DIA3
PIN DOA3
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER ME5 ;
  RECT 93.680 0.000 94.800 1.120 ;
  LAYER ME4 ;
  RECT 93.680 0.000 94.800 1.120 ;
  LAYER ME3 ;
  RECT 93.680 0.000 94.800 1.120 ;
  LAYER ME2 ;
  RECT 93.680 0.000 94.800 1.120 ;
  LAYER ME1 ;
  RECT 93.680 0.000 94.800 1.120 ;
 END
END DOA3
PIN DIA2
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER ME5 ;
  RECT 80.040 0.000 81.160 1.120 ;
  LAYER ME4 ;
  RECT 80.040 0.000 81.160 1.120 ;
  LAYER ME3 ;
  RECT 80.040 0.000 81.160 1.120 ;
  LAYER ME2 ;
  RECT 80.040 0.000 81.160 1.120 ;
  LAYER ME1 ;
  RECT 80.040 0.000 81.160 1.120 ;
 END
END DIA2
PIN DOA2
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME5 ;
  RECT 66.400 0.000 67.520 1.120 ;
  LAYER ME4 ;
  RECT 66.400 0.000 67.520 1.120 ;
  LAYER ME3 ;
  RECT 66.400 0.000 67.520 1.120 ;
  LAYER ME2 ;
  RECT 66.400 0.000 67.520 1.120 ;
  LAYER ME1 ;
  RECT 66.400 0.000 67.520 1.120 ;
 END
END DOA2
PIN DIA1
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER ME5 ;
  RECT 52.760 0.000 53.880 1.120 ;
  LAYER ME4 ;
  RECT 52.760 0.000 53.880 1.120 ;
  LAYER ME3 ;
  RECT 52.760 0.000 53.880 1.120 ;
  LAYER ME2 ;
  RECT 52.760 0.000 53.880 1.120 ;
  LAYER ME1 ;
  RECT 52.760 0.000 53.880 1.120 ;
 END
END DIA1
PIN DOA1
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME5 ;
  RECT 39.740 0.000 40.860 1.120 ;
  LAYER ME4 ;
  RECT 39.740 0.000 40.860 1.120 ;
  LAYER ME3 ;
  RECT 39.740 0.000 40.860 1.120 ;
  LAYER ME2 ;
  RECT 39.740 0.000 40.860 1.120 ;
  LAYER ME1 ;
  RECT 39.740 0.000 40.860 1.120 ;
 END
END DOA1
PIN DIA0
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER ME5 ;
  RECT 26.100 0.000 27.220 1.120 ;
  LAYER ME4 ;
  RECT 26.100 0.000 27.220 1.120 ;
  LAYER ME3 ;
  RECT 26.100 0.000 27.220 1.120 ;
  LAYER ME2 ;
  RECT 26.100 0.000 27.220 1.120 ;
  LAYER ME1 ;
  RECT 26.100 0.000 27.220 1.120 ;
 END
END DIA0
PIN DOA0
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER ME5 ;
  RECT 12.460 0.000 13.580 1.120 ;
  LAYER ME4 ;
  RECT 12.460 0.000 13.580 1.120 ;
  LAYER ME3 ;
  RECT 12.460 0.000 13.580 1.120 ;
  LAYER ME2 ;
  RECT 12.460 0.000 13.580 1.120 ;
  LAYER ME1 ;
  RECT 12.460 0.000 13.580 1.120 ;
 END
END DOA0
OBS
  LAYER ME1 SPACING 0.280 ;
  RECT 0.000 0.140 972.780 252.420 ;
  LAYER ME2 SPACING 0.320 ;
  RECT 0.000 0.140 972.780 252.420 ;
  LAYER ME3 SPACING 0.320 ;
  RECT 0.000 0.140 972.780 252.420 ;
  LAYER ME4 SPACING 0.600 ;
  RECT 0.000 0.140 972.780 252.420 ;
  LAYER VI1 ;
  RECT 0.000 0.140 972.780 252.420 ;
  LAYER VI2 ;
  RECT 0.000 0.140 972.780 252.420 ;
  LAYER VI3 ;
  RECT 0.000 0.140 972.780 252.420 ;
END
END DPSRAM_32_256
END LIBRARY



