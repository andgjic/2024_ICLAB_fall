# 
#              Synchronous High Speed Single Port SRAM Compiler 
# 
#                    UMC 0.18um GenericII Logic Process
#    __________________________________________________________________________
# 
# 
#      (C) Copyright 2002-2009 Faraday Technology Corp. All Rights Reserved.
#    
#    This source code is an unpublished work belongs to Faraday Technology
#    Corp.  It is considered a trade secret and is not to be divulged or
#    used by parties who have not received written authorization from
#    Faraday Technology Corp.
#    
#    Faraday's home page can be found at:
#    http://www.faraday-tech.com/
#   
#       Module Name      : Memory_32_256
#       Words            : 256
#       Bits             : 32
#       Byte-Write       : 1
#       Aspect Ratio     : 1
#       Output Loading   : 0.05  (pf)
#       Data Slew        : 0.02  (ns)
#       CK Slew          : 0.02  (ns)
#       Power Ring Width : 2  (um)
# 
# -----------------------------------------------------------------------------
# 
#       Library          : FSA0M_A
#       Memaker          : 200901.2.1
#       Date             : 2024/10/27 11:56:46
# 
# -----------------------------------------------------------------------------


NAMESCASESENSITIVE ON ;
MACRO Memory_32_256
CLASS BLOCK ;
FOREIGN Memory_32_256 0.000 0.000 ;
ORIGIN 0.000 0.000 ;
SIZE 542.500 BY 215.600 ;
SYMMETRY x y r90 ;
SITE core ;
PIN VCC
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
 PORT
  LAYER ME4 ;
  RECT 541.380 204.180 542.500 207.420 ;
  LAYER ME3 ;
  RECT 541.380 204.180 542.500 207.420 ;
  LAYER ME2 ;
  RECT 541.380 204.180 542.500 207.420 ;
  LAYER ME1 ;
  RECT 541.380 204.180 542.500 207.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 541.380 196.340 542.500 199.580 ;
  LAYER ME3 ;
  RECT 541.380 196.340 542.500 199.580 ;
  LAYER ME2 ;
  RECT 541.380 196.340 542.500 199.580 ;
  LAYER ME1 ;
  RECT 541.380 196.340 542.500 199.580 ;
 END
 PORT
  LAYER ME4 ;
  RECT 541.380 188.500 542.500 191.740 ;
  LAYER ME3 ;
  RECT 541.380 188.500 542.500 191.740 ;
  LAYER ME2 ;
  RECT 541.380 188.500 542.500 191.740 ;
  LAYER ME1 ;
  RECT 541.380 188.500 542.500 191.740 ;
 END
 PORT
  LAYER ME4 ;
  RECT 541.380 180.660 542.500 183.900 ;
  LAYER ME3 ;
  RECT 541.380 180.660 542.500 183.900 ;
  LAYER ME2 ;
  RECT 541.380 180.660 542.500 183.900 ;
  LAYER ME1 ;
  RECT 541.380 180.660 542.500 183.900 ;
 END
 PORT
  LAYER ME4 ;
  RECT 541.380 172.820 542.500 176.060 ;
  LAYER ME3 ;
  RECT 541.380 172.820 542.500 176.060 ;
  LAYER ME2 ;
  RECT 541.380 172.820 542.500 176.060 ;
  LAYER ME1 ;
  RECT 541.380 172.820 542.500 176.060 ;
 END
 PORT
  LAYER ME4 ;
  RECT 541.380 164.980 542.500 168.220 ;
  LAYER ME3 ;
  RECT 541.380 164.980 542.500 168.220 ;
  LAYER ME2 ;
  RECT 541.380 164.980 542.500 168.220 ;
  LAYER ME1 ;
  RECT 541.380 164.980 542.500 168.220 ;
 END
 PORT
  LAYER ME4 ;
  RECT 541.380 125.780 542.500 129.020 ;
  LAYER ME3 ;
  RECT 541.380 125.780 542.500 129.020 ;
  LAYER ME2 ;
  RECT 541.380 125.780 542.500 129.020 ;
  LAYER ME1 ;
  RECT 541.380 125.780 542.500 129.020 ;
 END
 PORT
  LAYER ME4 ;
  RECT 541.380 117.940 542.500 121.180 ;
  LAYER ME3 ;
  RECT 541.380 117.940 542.500 121.180 ;
  LAYER ME2 ;
  RECT 541.380 117.940 542.500 121.180 ;
  LAYER ME1 ;
  RECT 541.380 117.940 542.500 121.180 ;
 END
 PORT
  LAYER ME4 ;
  RECT 541.380 110.100 542.500 113.340 ;
  LAYER ME3 ;
  RECT 541.380 110.100 542.500 113.340 ;
  LAYER ME2 ;
  RECT 541.380 110.100 542.500 113.340 ;
  LAYER ME1 ;
  RECT 541.380 110.100 542.500 113.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 541.380 102.260 542.500 105.500 ;
  LAYER ME3 ;
  RECT 541.380 102.260 542.500 105.500 ;
  LAYER ME2 ;
  RECT 541.380 102.260 542.500 105.500 ;
  LAYER ME1 ;
  RECT 541.380 102.260 542.500 105.500 ;
 END
 PORT
  LAYER ME4 ;
  RECT 541.380 94.420 542.500 97.660 ;
  LAYER ME3 ;
  RECT 541.380 94.420 542.500 97.660 ;
  LAYER ME2 ;
  RECT 541.380 94.420 542.500 97.660 ;
  LAYER ME1 ;
  RECT 541.380 94.420 542.500 97.660 ;
 END
 PORT
  LAYER ME4 ;
  RECT 541.380 86.580 542.500 89.820 ;
  LAYER ME3 ;
  RECT 541.380 86.580 542.500 89.820 ;
  LAYER ME2 ;
  RECT 541.380 86.580 542.500 89.820 ;
  LAYER ME1 ;
  RECT 541.380 86.580 542.500 89.820 ;
 END
 PORT
  LAYER ME4 ;
  RECT 541.380 47.380 542.500 50.620 ;
  LAYER ME3 ;
  RECT 541.380 47.380 542.500 50.620 ;
  LAYER ME2 ;
  RECT 541.380 47.380 542.500 50.620 ;
  LAYER ME1 ;
  RECT 541.380 47.380 542.500 50.620 ;
 END
 PORT
  LAYER ME4 ;
  RECT 541.380 39.540 542.500 42.780 ;
  LAYER ME3 ;
  RECT 541.380 39.540 542.500 42.780 ;
  LAYER ME2 ;
  RECT 541.380 39.540 542.500 42.780 ;
  LAYER ME1 ;
  RECT 541.380 39.540 542.500 42.780 ;
 END
 PORT
  LAYER ME4 ;
  RECT 541.380 31.700 542.500 34.940 ;
  LAYER ME3 ;
  RECT 541.380 31.700 542.500 34.940 ;
  LAYER ME2 ;
  RECT 541.380 31.700 542.500 34.940 ;
  LAYER ME1 ;
  RECT 541.380 31.700 542.500 34.940 ;
 END
 PORT
  LAYER ME4 ;
  RECT 541.380 23.860 542.500 27.100 ;
  LAYER ME3 ;
  RECT 541.380 23.860 542.500 27.100 ;
  LAYER ME2 ;
  RECT 541.380 23.860 542.500 27.100 ;
  LAYER ME1 ;
  RECT 541.380 23.860 542.500 27.100 ;
 END
 PORT
  LAYER ME4 ;
  RECT 541.380 16.020 542.500 19.260 ;
  LAYER ME3 ;
  RECT 541.380 16.020 542.500 19.260 ;
  LAYER ME2 ;
  RECT 541.380 16.020 542.500 19.260 ;
  LAYER ME1 ;
  RECT 541.380 16.020 542.500 19.260 ;
 END
 PORT
  LAYER ME4 ;
  RECT 541.380 8.180 542.500 11.420 ;
  LAYER ME3 ;
  RECT 541.380 8.180 542.500 11.420 ;
  LAYER ME2 ;
  RECT 541.380 8.180 542.500 11.420 ;
  LAYER ME1 ;
  RECT 541.380 8.180 542.500 11.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 204.180 1.120 207.420 ;
  LAYER ME3 ;
  RECT 0.000 204.180 1.120 207.420 ;
  LAYER ME2 ;
  RECT 0.000 204.180 1.120 207.420 ;
  LAYER ME1 ;
  RECT 0.000 204.180 1.120 207.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 196.340 1.120 199.580 ;
  LAYER ME3 ;
  RECT 0.000 196.340 1.120 199.580 ;
  LAYER ME2 ;
  RECT 0.000 196.340 1.120 199.580 ;
  LAYER ME1 ;
  RECT 0.000 196.340 1.120 199.580 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 188.500 1.120 191.740 ;
  LAYER ME3 ;
  RECT 0.000 188.500 1.120 191.740 ;
  LAYER ME2 ;
  RECT 0.000 188.500 1.120 191.740 ;
  LAYER ME1 ;
  RECT 0.000 188.500 1.120 191.740 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 180.660 1.120 183.900 ;
  LAYER ME3 ;
  RECT 0.000 180.660 1.120 183.900 ;
  LAYER ME2 ;
  RECT 0.000 180.660 1.120 183.900 ;
  LAYER ME1 ;
  RECT 0.000 180.660 1.120 183.900 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 172.820 1.120 176.060 ;
  LAYER ME3 ;
  RECT 0.000 172.820 1.120 176.060 ;
  LAYER ME2 ;
  RECT 0.000 172.820 1.120 176.060 ;
  LAYER ME1 ;
  RECT 0.000 172.820 1.120 176.060 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 164.980 1.120 168.220 ;
  LAYER ME3 ;
  RECT 0.000 164.980 1.120 168.220 ;
  LAYER ME2 ;
  RECT 0.000 164.980 1.120 168.220 ;
  LAYER ME1 ;
  RECT 0.000 164.980 1.120 168.220 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 125.780 1.120 129.020 ;
  LAYER ME3 ;
  RECT 0.000 125.780 1.120 129.020 ;
  LAYER ME2 ;
  RECT 0.000 125.780 1.120 129.020 ;
  LAYER ME1 ;
  RECT 0.000 125.780 1.120 129.020 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 117.940 1.120 121.180 ;
  LAYER ME3 ;
  RECT 0.000 117.940 1.120 121.180 ;
  LAYER ME2 ;
  RECT 0.000 117.940 1.120 121.180 ;
  LAYER ME1 ;
  RECT 0.000 117.940 1.120 121.180 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 110.100 1.120 113.340 ;
  LAYER ME3 ;
  RECT 0.000 110.100 1.120 113.340 ;
  LAYER ME2 ;
  RECT 0.000 110.100 1.120 113.340 ;
  LAYER ME1 ;
  RECT 0.000 110.100 1.120 113.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 102.260 1.120 105.500 ;
  LAYER ME3 ;
  RECT 0.000 102.260 1.120 105.500 ;
  LAYER ME2 ;
  RECT 0.000 102.260 1.120 105.500 ;
  LAYER ME1 ;
  RECT 0.000 102.260 1.120 105.500 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 94.420 1.120 97.660 ;
  LAYER ME3 ;
  RECT 0.000 94.420 1.120 97.660 ;
  LAYER ME2 ;
  RECT 0.000 94.420 1.120 97.660 ;
  LAYER ME1 ;
  RECT 0.000 94.420 1.120 97.660 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 86.580 1.120 89.820 ;
  LAYER ME3 ;
  RECT 0.000 86.580 1.120 89.820 ;
  LAYER ME2 ;
  RECT 0.000 86.580 1.120 89.820 ;
  LAYER ME1 ;
  RECT 0.000 86.580 1.120 89.820 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 47.380 1.120 50.620 ;
  LAYER ME3 ;
  RECT 0.000 47.380 1.120 50.620 ;
  LAYER ME2 ;
  RECT 0.000 47.380 1.120 50.620 ;
  LAYER ME1 ;
  RECT 0.000 47.380 1.120 50.620 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 39.540 1.120 42.780 ;
  LAYER ME3 ;
  RECT 0.000 39.540 1.120 42.780 ;
  LAYER ME2 ;
  RECT 0.000 39.540 1.120 42.780 ;
  LAYER ME1 ;
  RECT 0.000 39.540 1.120 42.780 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 31.700 1.120 34.940 ;
  LAYER ME3 ;
  RECT 0.000 31.700 1.120 34.940 ;
  LAYER ME2 ;
  RECT 0.000 31.700 1.120 34.940 ;
  LAYER ME1 ;
  RECT 0.000 31.700 1.120 34.940 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 23.860 1.120 27.100 ;
  LAYER ME3 ;
  RECT 0.000 23.860 1.120 27.100 ;
  LAYER ME2 ;
  RECT 0.000 23.860 1.120 27.100 ;
  LAYER ME1 ;
  RECT 0.000 23.860 1.120 27.100 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 16.020 1.120 19.260 ;
  LAYER ME3 ;
  RECT 0.000 16.020 1.120 19.260 ;
  LAYER ME2 ;
  RECT 0.000 16.020 1.120 19.260 ;
  LAYER ME1 ;
  RECT 0.000 16.020 1.120 19.260 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 8.180 1.120 11.420 ;
  LAYER ME3 ;
  RECT 0.000 8.180 1.120 11.420 ;
  LAYER ME2 ;
  RECT 0.000 8.180 1.120 11.420 ;
  LAYER ME1 ;
  RECT 0.000 8.180 1.120 11.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 528.640 214.480 532.180 215.600 ;
  LAYER ME3 ;
  RECT 528.640 214.480 532.180 215.600 ;
  LAYER ME2 ;
  RECT 528.640 214.480 532.180 215.600 ;
  LAYER ME1 ;
  RECT 528.640 214.480 532.180 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 485.240 214.480 488.780 215.600 ;
  LAYER ME3 ;
  RECT 485.240 214.480 488.780 215.600 ;
  LAYER ME2 ;
  RECT 485.240 214.480 488.780 215.600 ;
  LAYER ME1 ;
  RECT 485.240 214.480 488.780 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 476.560 214.480 480.100 215.600 ;
  LAYER ME3 ;
  RECT 476.560 214.480 480.100 215.600 ;
  LAYER ME2 ;
  RECT 476.560 214.480 480.100 215.600 ;
  LAYER ME1 ;
  RECT 476.560 214.480 480.100 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 467.880 214.480 471.420 215.600 ;
  LAYER ME3 ;
  RECT 467.880 214.480 471.420 215.600 ;
  LAYER ME2 ;
  RECT 467.880 214.480 471.420 215.600 ;
  LAYER ME1 ;
  RECT 467.880 214.480 471.420 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 459.200 214.480 462.740 215.600 ;
  LAYER ME3 ;
  RECT 459.200 214.480 462.740 215.600 ;
  LAYER ME2 ;
  RECT 459.200 214.480 462.740 215.600 ;
  LAYER ME1 ;
  RECT 459.200 214.480 462.740 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 450.520 214.480 454.060 215.600 ;
  LAYER ME3 ;
  RECT 450.520 214.480 454.060 215.600 ;
  LAYER ME2 ;
  RECT 450.520 214.480 454.060 215.600 ;
  LAYER ME1 ;
  RECT 450.520 214.480 454.060 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 441.840 214.480 445.380 215.600 ;
  LAYER ME3 ;
  RECT 441.840 214.480 445.380 215.600 ;
  LAYER ME2 ;
  RECT 441.840 214.480 445.380 215.600 ;
  LAYER ME1 ;
  RECT 441.840 214.480 445.380 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 398.440 214.480 401.980 215.600 ;
  LAYER ME3 ;
  RECT 398.440 214.480 401.980 215.600 ;
  LAYER ME2 ;
  RECT 398.440 214.480 401.980 215.600 ;
  LAYER ME1 ;
  RECT 398.440 214.480 401.980 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 389.760 214.480 393.300 215.600 ;
  LAYER ME3 ;
  RECT 389.760 214.480 393.300 215.600 ;
  LAYER ME2 ;
  RECT 389.760 214.480 393.300 215.600 ;
  LAYER ME1 ;
  RECT 389.760 214.480 393.300 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 381.080 214.480 384.620 215.600 ;
  LAYER ME3 ;
  RECT 381.080 214.480 384.620 215.600 ;
  LAYER ME2 ;
  RECT 381.080 214.480 384.620 215.600 ;
  LAYER ME1 ;
  RECT 381.080 214.480 384.620 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 372.400 214.480 375.940 215.600 ;
  LAYER ME3 ;
  RECT 372.400 214.480 375.940 215.600 ;
  LAYER ME2 ;
  RECT 372.400 214.480 375.940 215.600 ;
  LAYER ME1 ;
  RECT 372.400 214.480 375.940 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 363.720 214.480 367.260 215.600 ;
  LAYER ME3 ;
  RECT 363.720 214.480 367.260 215.600 ;
  LAYER ME2 ;
  RECT 363.720 214.480 367.260 215.600 ;
  LAYER ME1 ;
  RECT 363.720 214.480 367.260 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 355.040 214.480 358.580 215.600 ;
  LAYER ME3 ;
  RECT 355.040 214.480 358.580 215.600 ;
  LAYER ME2 ;
  RECT 355.040 214.480 358.580 215.600 ;
  LAYER ME1 ;
  RECT 355.040 214.480 358.580 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 311.640 214.480 315.180 215.600 ;
  LAYER ME3 ;
  RECT 311.640 214.480 315.180 215.600 ;
  LAYER ME2 ;
  RECT 311.640 214.480 315.180 215.600 ;
  LAYER ME1 ;
  RECT 311.640 214.480 315.180 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 302.960 214.480 306.500 215.600 ;
  LAYER ME3 ;
  RECT 302.960 214.480 306.500 215.600 ;
  LAYER ME2 ;
  RECT 302.960 214.480 306.500 215.600 ;
  LAYER ME1 ;
  RECT 302.960 214.480 306.500 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 294.280 214.480 297.820 215.600 ;
  LAYER ME3 ;
  RECT 294.280 214.480 297.820 215.600 ;
  LAYER ME2 ;
  RECT 294.280 214.480 297.820 215.600 ;
  LAYER ME1 ;
  RECT 294.280 214.480 297.820 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 285.600 214.480 289.140 215.600 ;
  LAYER ME3 ;
  RECT 285.600 214.480 289.140 215.600 ;
  LAYER ME2 ;
  RECT 285.600 214.480 289.140 215.600 ;
  LAYER ME1 ;
  RECT 285.600 214.480 289.140 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 276.920 214.480 280.460 215.600 ;
  LAYER ME3 ;
  RECT 276.920 214.480 280.460 215.600 ;
  LAYER ME2 ;
  RECT 276.920 214.480 280.460 215.600 ;
  LAYER ME1 ;
  RECT 276.920 214.480 280.460 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 268.240 214.480 271.780 215.600 ;
  LAYER ME3 ;
  RECT 268.240 214.480 271.780 215.600 ;
  LAYER ME2 ;
  RECT 268.240 214.480 271.780 215.600 ;
  LAYER ME1 ;
  RECT 268.240 214.480 271.780 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 224.840 214.480 228.380 215.600 ;
  LAYER ME3 ;
  RECT 224.840 214.480 228.380 215.600 ;
  LAYER ME2 ;
  RECT 224.840 214.480 228.380 215.600 ;
  LAYER ME1 ;
  RECT 224.840 214.480 228.380 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 216.160 214.480 219.700 215.600 ;
  LAYER ME3 ;
  RECT 216.160 214.480 219.700 215.600 ;
  LAYER ME2 ;
  RECT 216.160 214.480 219.700 215.600 ;
  LAYER ME1 ;
  RECT 216.160 214.480 219.700 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 207.480 214.480 211.020 215.600 ;
  LAYER ME3 ;
  RECT 207.480 214.480 211.020 215.600 ;
  LAYER ME2 ;
  RECT 207.480 214.480 211.020 215.600 ;
  LAYER ME1 ;
  RECT 207.480 214.480 211.020 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 198.800 214.480 202.340 215.600 ;
  LAYER ME3 ;
  RECT 198.800 214.480 202.340 215.600 ;
  LAYER ME2 ;
  RECT 198.800 214.480 202.340 215.600 ;
  LAYER ME1 ;
  RECT 198.800 214.480 202.340 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 190.120 214.480 193.660 215.600 ;
  LAYER ME3 ;
  RECT 190.120 214.480 193.660 215.600 ;
  LAYER ME2 ;
  RECT 190.120 214.480 193.660 215.600 ;
  LAYER ME1 ;
  RECT 190.120 214.480 193.660 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 181.440 214.480 184.980 215.600 ;
  LAYER ME3 ;
  RECT 181.440 214.480 184.980 215.600 ;
  LAYER ME2 ;
  RECT 181.440 214.480 184.980 215.600 ;
  LAYER ME1 ;
  RECT 181.440 214.480 184.980 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 138.040 214.480 141.580 215.600 ;
  LAYER ME3 ;
  RECT 138.040 214.480 141.580 215.600 ;
  LAYER ME2 ;
  RECT 138.040 214.480 141.580 215.600 ;
  LAYER ME1 ;
  RECT 138.040 214.480 141.580 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 129.360 214.480 132.900 215.600 ;
  LAYER ME3 ;
  RECT 129.360 214.480 132.900 215.600 ;
  LAYER ME2 ;
  RECT 129.360 214.480 132.900 215.600 ;
  LAYER ME1 ;
  RECT 129.360 214.480 132.900 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 120.680 214.480 124.220 215.600 ;
  LAYER ME3 ;
  RECT 120.680 214.480 124.220 215.600 ;
  LAYER ME2 ;
  RECT 120.680 214.480 124.220 215.600 ;
  LAYER ME1 ;
  RECT 120.680 214.480 124.220 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 112.000 214.480 115.540 215.600 ;
  LAYER ME3 ;
  RECT 112.000 214.480 115.540 215.600 ;
  LAYER ME2 ;
  RECT 112.000 214.480 115.540 215.600 ;
  LAYER ME1 ;
  RECT 112.000 214.480 115.540 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 103.320 214.480 106.860 215.600 ;
  LAYER ME3 ;
  RECT 103.320 214.480 106.860 215.600 ;
  LAYER ME2 ;
  RECT 103.320 214.480 106.860 215.600 ;
  LAYER ME1 ;
  RECT 103.320 214.480 106.860 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 94.640 214.480 98.180 215.600 ;
  LAYER ME3 ;
  RECT 94.640 214.480 98.180 215.600 ;
  LAYER ME2 ;
  RECT 94.640 214.480 98.180 215.600 ;
  LAYER ME1 ;
  RECT 94.640 214.480 98.180 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 51.240 214.480 54.780 215.600 ;
  LAYER ME3 ;
  RECT 51.240 214.480 54.780 215.600 ;
  LAYER ME2 ;
  RECT 51.240 214.480 54.780 215.600 ;
  LAYER ME1 ;
  RECT 51.240 214.480 54.780 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 42.560 214.480 46.100 215.600 ;
  LAYER ME3 ;
  RECT 42.560 214.480 46.100 215.600 ;
  LAYER ME2 ;
  RECT 42.560 214.480 46.100 215.600 ;
  LAYER ME1 ;
  RECT 42.560 214.480 46.100 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 33.880 214.480 37.420 215.600 ;
  LAYER ME3 ;
  RECT 33.880 214.480 37.420 215.600 ;
  LAYER ME2 ;
  RECT 33.880 214.480 37.420 215.600 ;
  LAYER ME1 ;
  RECT 33.880 214.480 37.420 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 25.200 214.480 28.740 215.600 ;
  LAYER ME3 ;
  RECT 25.200 214.480 28.740 215.600 ;
  LAYER ME2 ;
  RECT 25.200 214.480 28.740 215.600 ;
  LAYER ME1 ;
  RECT 25.200 214.480 28.740 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 16.520 214.480 20.060 215.600 ;
  LAYER ME3 ;
  RECT 16.520 214.480 20.060 215.600 ;
  LAYER ME2 ;
  RECT 16.520 214.480 20.060 215.600 ;
  LAYER ME1 ;
  RECT 16.520 214.480 20.060 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 7.840 214.480 11.380 215.600 ;
  LAYER ME3 ;
  RECT 7.840 214.480 11.380 215.600 ;
  LAYER ME2 ;
  RECT 7.840 214.480 11.380 215.600 ;
  LAYER ME1 ;
  RECT 7.840 214.480 11.380 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 522.440 0.000 525.980 1.120 ;
  LAYER ME3 ;
  RECT 522.440 0.000 525.980 1.120 ;
  LAYER ME2 ;
  RECT 522.440 0.000 525.980 1.120 ;
  LAYER ME1 ;
  RECT 522.440 0.000 525.980 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 500.740 0.000 504.280 1.120 ;
  LAYER ME3 ;
  RECT 500.740 0.000 504.280 1.120 ;
  LAYER ME2 ;
  RECT 500.740 0.000 504.280 1.120 ;
  LAYER ME1 ;
  RECT 500.740 0.000 504.280 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 479.660 0.000 483.200 1.120 ;
  LAYER ME3 ;
  RECT 479.660 0.000 483.200 1.120 ;
  LAYER ME2 ;
  RECT 479.660 0.000 483.200 1.120 ;
  LAYER ME1 ;
  RECT 479.660 0.000 483.200 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 453.000 0.000 456.540 1.120 ;
  LAYER ME3 ;
  RECT 453.000 0.000 456.540 1.120 ;
  LAYER ME2 ;
  RECT 453.000 0.000 456.540 1.120 ;
  LAYER ME1 ;
  RECT 453.000 0.000 456.540 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 339.540 0.000 343.080 1.120 ;
  LAYER ME3 ;
  RECT 339.540 0.000 343.080 1.120 ;
  LAYER ME2 ;
  RECT 339.540 0.000 343.080 1.120 ;
  LAYER ME1 ;
  RECT 339.540 0.000 343.080 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 322.800 0.000 326.340 1.120 ;
  LAYER ME3 ;
  RECT 322.800 0.000 326.340 1.120 ;
  LAYER ME2 ;
  RECT 322.800 0.000 326.340 1.120 ;
  LAYER ME1 ;
  RECT 322.800 0.000 326.340 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 286.840 0.000 290.380 1.120 ;
  LAYER ME3 ;
  RECT 286.840 0.000 290.380 1.120 ;
  LAYER ME2 ;
  RECT 286.840 0.000 290.380 1.120 ;
  LAYER ME1 ;
  RECT 286.840 0.000 290.380 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 278.160 0.000 281.700 1.120 ;
  LAYER ME3 ;
  RECT 278.160 0.000 281.700 1.120 ;
  LAYER ME2 ;
  RECT 278.160 0.000 281.700 1.120 ;
  LAYER ME1 ;
  RECT 278.160 0.000 281.700 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 257.080 0.000 260.620 1.120 ;
  LAYER ME3 ;
  RECT 257.080 0.000 260.620 1.120 ;
  LAYER ME2 ;
  RECT 257.080 0.000 260.620 1.120 ;
  LAYER ME1 ;
  RECT 257.080 0.000 260.620 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 235.380 0.000 238.920 1.120 ;
  LAYER ME3 ;
  RECT 235.380 0.000 238.920 1.120 ;
  LAYER ME2 ;
  RECT 235.380 0.000 238.920 1.120 ;
  LAYER ME1 ;
  RECT 235.380 0.000 238.920 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 126.880 0.000 130.420 1.120 ;
  LAYER ME3 ;
  RECT 126.880 0.000 130.420 1.120 ;
  LAYER ME2 ;
  RECT 126.880 0.000 130.420 1.120 ;
  LAYER ME1 ;
  RECT 126.880 0.000 130.420 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 100.220 0.000 103.760 1.120 ;
  LAYER ME3 ;
  RECT 100.220 0.000 103.760 1.120 ;
  LAYER ME2 ;
  RECT 100.220 0.000 103.760 1.120 ;
  LAYER ME1 ;
  RECT 100.220 0.000 103.760 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 83.480 0.000 87.020 1.120 ;
  LAYER ME3 ;
  RECT 83.480 0.000 87.020 1.120 ;
  LAYER ME2 ;
  RECT 83.480 0.000 87.020 1.120 ;
  LAYER ME1 ;
  RECT 83.480 0.000 87.020 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 56.820 0.000 60.360 1.120 ;
  LAYER ME3 ;
  RECT 56.820 0.000 60.360 1.120 ;
  LAYER ME2 ;
  RECT 56.820 0.000 60.360 1.120 ;
  LAYER ME1 ;
  RECT 56.820 0.000 60.360 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 35.740 0.000 39.280 1.120 ;
  LAYER ME3 ;
  RECT 35.740 0.000 39.280 1.120 ;
  LAYER ME2 ;
  RECT 35.740 0.000 39.280 1.120 ;
  LAYER ME1 ;
  RECT 35.740 0.000 39.280 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 14.040 0.000 17.580 1.120 ;
  LAYER ME3 ;
  RECT 14.040 0.000 17.580 1.120 ;
  LAYER ME2 ;
  RECT 14.040 0.000 17.580 1.120 ;
  LAYER ME1 ;
  RECT 14.040 0.000 17.580 1.120 ;
 END
END VCC
PIN GND
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
 PORT
  LAYER ME4 ;
  RECT 541.380 200.260 542.500 203.500 ;
  LAYER ME3 ;
  RECT 541.380 200.260 542.500 203.500 ;
  LAYER ME2 ;
  RECT 541.380 200.260 542.500 203.500 ;
  LAYER ME1 ;
  RECT 541.380 200.260 542.500 203.500 ;
 END
 PORT
  LAYER ME4 ;
  RECT 541.380 192.420 542.500 195.660 ;
  LAYER ME3 ;
  RECT 541.380 192.420 542.500 195.660 ;
  LAYER ME2 ;
  RECT 541.380 192.420 542.500 195.660 ;
  LAYER ME1 ;
  RECT 541.380 192.420 542.500 195.660 ;
 END
 PORT
  LAYER ME4 ;
  RECT 541.380 184.580 542.500 187.820 ;
  LAYER ME3 ;
  RECT 541.380 184.580 542.500 187.820 ;
  LAYER ME2 ;
  RECT 541.380 184.580 542.500 187.820 ;
  LAYER ME1 ;
  RECT 541.380 184.580 542.500 187.820 ;
 END
 PORT
  LAYER ME4 ;
  RECT 541.380 176.740 542.500 179.980 ;
  LAYER ME3 ;
  RECT 541.380 176.740 542.500 179.980 ;
  LAYER ME2 ;
  RECT 541.380 176.740 542.500 179.980 ;
  LAYER ME1 ;
  RECT 541.380 176.740 542.500 179.980 ;
 END
 PORT
  LAYER ME4 ;
  RECT 541.380 168.900 542.500 172.140 ;
  LAYER ME3 ;
  RECT 541.380 168.900 542.500 172.140 ;
  LAYER ME2 ;
  RECT 541.380 168.900 542.500 172.140 ;
  LAYER ME1 ;
  RECT 541.380 168.900 542.500 172.140 ;
 END
 PORT
  LAYER ME4 ;
  RECT 541.380 129.700 542.500 132.940 ;
  LAYER ME3 ;
  RECT 541.380 129.700 542.500 132.940 ;
  LAYER ME2 ;
  RECT 541.380 129.700 542.500 132.940 ;
  LAYER ME1 ;
  RECT 541.380 129.700 542.500 132.940 ;
 END
 PORT
  LAYER ME4 ;
  RECT 541.380 121.860 542.500 125.100 ;
  LAYER ME3 ;
  RECT 541.380 121.860 542.500 125.100 ;
  LAYER ME2 ;
  RECT 541.380 121.860 542.500 125.100 ;
  LAYER ME1 ;
  RECT 541.380 121.860 542.500 125.100 ;
 END
 PORT
  LAYER ME4 ;
  RECT 541.380 114.020 542.500 117.260 ;
  LAYER ME3 ;
  RECT 541.380 114.020 542.500 117.260 ;
  LAYER ME2 ;
  RECT 541.380 114.020 542.500 117.260 ;
  LAYER ME1 ;
  RECT 541.380 114.020 542.500 117.260 ;
 END
 PORT
  LAYER ME4 ;
  RECT 541.380 106.180 542.500 109.420 ;
  LAYER ME3 ;
  RECT 541.380 106.180 542.500 109.420 ;
  LAYER ME2 ;
  RECT 541.380 106.180 542.500 109.420 ;
  LAYER ME1 ;
  RECT 541.380 106.180 542.500 109.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 541.380 98.340 542.500 101.580 ;
  LAYER ME3 ;
  RECT 541.380 98.340 542.500 101.580 ;
  LAYER ME2 ;
  RECT 541.380 98.340 542.500 101.580 ;
  LAYER ME1 ;
  RECT 541.380 98.340 542.500 101.580 ;
 END
 PORT
  LAYER ME4 ;
  RECT 541.380 90.500 542.500 93.740 ;
  LAYER ME3 ;
  RECT 541.380 90.500 542.500 93.740 ;
  LAYER ME2 ;
  RECT 541.380 90.500 542.500 93.740 ;
  LAYER ME1 ;
  RECT 541.380 90.500 542.500 93.740 ;
 END
 PORT
  LAYER ME4 ;
  RECT 541.380 51.300 542.500 54.540 ;
  LAYER ME3 ;
  RECT 541.380 51.300 542.500 54.540 ;
  LAYER ME2 ;
  RECT 541.380 51.300 542.500 54.540 ;
  LAYER ME1 ;
  RECT 541.380 51.300 542.500 54.540 ;
 END
 PORT
  LAYER ME4 ;
  RECT 541.380 43.460 542.500 46.700 ;
  LAYER ME3 ;
  RECT 541.380 43.460 542.500 46.700 ;
  LAYER ME2 ;
  RECT 541.380 43.460 542.500 46.700 ;
  LAYER ME1 ;
  RECT 541.380 43.460 542.500 46.700 ;
 END
 PORT
  LAYER ME4 ;
  RECT 541.380 35.620 542.500 38.860 ;
  LAYER ME3 ;
  RECT 541.380 35.620 542.500 38.860 ;
  LAYER ME2 ;
  RECT 541.380 35.620 542.500 38.860 ;
  LAYER ME1 ;
  RECT 541.380 35.620 542.500 38.860 ;
 END
 PORT
  LAYER ME4 ;
  RECT 541.380 27.780 542.500 31.020 ;
  LAYER ME3 ;
  RECT 541.380 27.780 542.500 31.020 ;
  LAYER ME2 ;
  RECT 541.380 27.780 542.500 31.020 ;
  LAYER ME1 ;
  RECT 541.380 27.780 542.500 31.020 ;
 END
 PORT
  LAYER ME4 ;
  RECT 541.380 19.940 542.500 23.180 ;
  LAYER ME3 ;
  RECT 541.380 19.940 542.500 23.180 ;
  LAYER ME2 ;
  RECT 541.380 19.940 542.500 23.180 ;
  LAYER ME1 ;
  RECT 541.380 19.940 542.500 23.180 ;
 END
 PORT
  LAYER ME4 ;
  RECT 541.380 12.100 542.500 15.340 ;
  LAYER ME3 ;
  RECT 541.380 12.100 542.500 15.340 ;
  LAYER ME2 ;
  RECT 541.380 12.100 542.500 15.340 ;
  LAYER ME1 ;
  RECT 541.380 12.100 542.500 15.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 200.260 1.120 203.500 ;
  LAYER ME3 ;
  RECT 0.000 200.260 1.120 203.500 ;
  LAYER ME2 ;
  RECT 0.000 200.260 1.120 203.500 ;
  LAYER ME1 ;
  RECT 0.000 200.260 1.120 203.500 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 192.420 1.120 195.660 ;
  LAYER ME3 ;
  RECT 0.000 192.420 1.120 195.660 ;
  LAYER ME2 ;
  RECT 0.000 192.420 1.120 195.660 ;
  LAYER ME1 ;
  RECT 0.000 192.420 1.120 195.660 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 184.580 1.120 187.820 ;
  LAYER ME3 ;
  RECT 0.000 184.580 1.120 187.820 ;
  LAYER ME2 ;
  RECT 0.000 184.580 1.120 187.820 ;
  LAYER ME1 ;
  RECT 0.000 184.580 1.120 187.820 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 176.740 1.120 179.980 ;
  LAYER ME3 ;
  RECT 0.000 176.740 1.120 179.980 ;
  LAYER ME2 ;
  RECT 0.000 176.740 1.120 179.980 ;
  LAYER ME1 ;
  RECT 0.000 176.740 1.120 179.980 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 168.900 1.120 172.140 ;
  LAYER ME3 ;
  RECT 0.000 168.900 1.120 172.140 ;
  LAYER ME2 ;
  RECT 0.000 168.900 1.120 172.140 ;
  LAYER ME1 ;
  RECT 0.000 168.900 1.120 172.140 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 129.700 1.120 132.940 ;
  LAYER ME3 ;
  RECT 0.000 129.700 1.120 132.940 ;
  LAYER ME2 ;
  RECT 0.000 129.700 1.120 132.940 ;
  LAYER ME1 ;
  RECT 0.000 129.700 1.120 132.940 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 121.860 1.120 125.100 ;
  LAYER ME3 ;
  RECT 0.000 121.860 1.120 125.100 ;
  LAYER ME2 ;
  RECT 0.000 121.860 1.120 125.100 ;
  LAYER ME1 ;
  RECT 0.000 121.860 1.120 125.100 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 114.020 1.120 117.260 ;
  LAYER ME3 ;
  RECT 0.000 114.020 1.120 117.260 ;
  LAYER ME2 ;
  RECT 0.000 114.020 1.120 117.260 ;
  LAYER ME1 ;
  RECT 0.000 114.020 1.120 117.260 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 106.180 1.120 109.420 ;
  LAYER ME3 ;
  RECT 0.000 106.180 1.120 109.420 ;
  LAYER ME2 ;
  RECT 0.000 106.180 1.120 109.420 ;
  LAYER ME1 ;
  RECT 0.000 106.180 1.120 109.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 98.340 1.120 101.580 ;
  LAYER ME3 ;
  RECT 0.000 98.340 1.120 101.580 ;
  LAYER ME2 ;
  RECT 0.000 98.340 1.120 101.580 ;
  LAYER ME1 ;
  RECT 0.000 98.340 1.120 101.580 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 90.500 1.120 93.740 ;
  LAYER ME3 ;
  RECT 0.000 90.500 1.120 93.740 ;
  LAYER ME2 ;
  RECT 0.000 90.500 1.120 93.740 ;
  LAYER ME1 ;
  RECT 0.000 90.500 1.120 93.740 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 51.300 1.120 54.540 ;
  LAYER ME3 ;
  RECT 0.000 51.300 1.120 54.540 ;
  LAYER ME2 ;
  RECT 0.000 51.300 1.120 54.540 ;
  LAYER ME1 ;
  RECT 0.000 51.300 1.120 54.540 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 43.460 1.120 46.700 ;
  LAYER ME3 ;
  RECT 0.000 43.460 1.120 46.700 ;
  LAYER ME2 ;
  RECT 0.000 43.460 1.120 46.700 ;
  LAYER ME1 ;
  RECT 0.000 43.460 1.120 46.700 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 35.620 1.120 38.860 ;
  LAYER ME3 ;
  RECT 0.000 35.620 1.120 38.860 ;
  LAYER ME2 ;
  RECT 0.000 35.620 1.120 38.860 ;
  LAYER ME1 ;
  RECT 0.000 35.620 1.120 38.860 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 27.780 1.120 31.020 ;
  LAYER ME3 ;
  RECT 0.000 27.780 1.120 31.020 ;
  LAYER ME2 ;
  RECT 0.000 27.780 1.120 31.020 ;
  LAYER ME1 ;
  RECT 0.000 27.780 1.120 31.020 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 19.940 1.120 23.180 ;
  LAYER ME3 ;
  RECT 0.000 19.940 1.120 23.180 ;
  LAYER ME2 ;
  RECT 0.000 19.940 1.120 23.180 ;
  LAYER ME1 ;
  RECT 0.000 19.940 1.120 23.180 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 12.100 1.120 15.340 ;
  LAYER ME3 ;
  RECT 0.000 12.100 1.120 15.340 ;
  LAYER ME2 ;
  RECT 0.000 12.100 1.120 15.340 ;
  LAYER ME1 ;
  RECT 0.000 12.100 1.120 15.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 489.580 214.480 493.120 215.600 ;
  LAYER ME3 ;
  RECT 489.580 214.480 493.120 215.600 ;
  LAYER ME2 ;
  RECT 489.580 214.480 493.120 215.600 ;
  LAYER ME1 ;
  RECT 489.580 214.480 493.120 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 480.900 214.480 484.440 215.600 ;
  LAYER ME3 ;
  RECT 480.900 214.480 484.440 215.600 ;
  LAYER ME2 ;
  RECT 480.900 214.480 484.440 215.600 ;
  LAYER ME1 ;
  RECT 480.900 214.480 484.440 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 472.220 214.480 475.760 215.600 ;
  LAYER ME3 ;
  RECT 472.220 214.480 475.760 215.600 ;
  LAYER ME2 ;
  RECT 472.220 214.480 475.760 215.600 ;
  LAYER ME1 ;
  RECT 472.220 214.480 475.760 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 463.540 214.480 467.080 215.600 ;
  LAYER ME3 ;
  RECT 463.540 214.480 467.080 215.600 ;
  LAYER ME2 ;
  RECT 463.540 214.480 467.080 215.600 ;
  LAYER ME1 ;
  RECT 463.540 214.480 467.080 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 454.860 214.480 458.400 215.600 ;
  LAYER ME3 ;
  RECT 454.860 214.480 458.400 215.600 ;
  LAYER ME2 ;
  RECT 454.860 214.480 458.400 215.600 ;
  LAYER ME1 ;
  RECT 454.860 214.480 458.400 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 446.180 214.480 449.720 215.600 ;
  LAYER ME3 ;
  RECT 446.180 214.480 449.720 215.600 ;
  LAYER ME2 ;
  RECT 446.180 214.480 449.720 215.600 ;
  LAYER ME1 ;
  RECT 446.180 214.480 449.720 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 402.780 214.480 406.320 215.600 ;
  LAYER ME3 ;
  RECT 402.780 214.480 406.320 215.600 ;
  LAYER ME2 ;
  RECT 402.780 214.480 406.320 215.600 ;
  LAYER ME1 ;
  RECT 402.780 214.480 406.320 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 394.100 214.480 397.640 215.600 ;
  LAYER ME3 ;
  RECT 394.100 214.480 397.640 215.600 ;
  LAYER ME2 ;
  RECT 394.100 214.480 397.640 215.600 ;
  LAYER ME1 ;
  RECT 394.100 214.480 397.640 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 385.420 214.480 388.960 215.600 ;
  LAYER ME3 ;
  RECT 385.420 214.480 388.960 215.600 ;
  LAYER ME2 ;
  RECT 385.420 214.480 388.960 215.600 ;
  LAYER ME1 ;
  RECT 385.420 214.480 388.960 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 376.740 214.480 380.280 215.600 ;
  LAYER ME3 ;
  RECT 376.740 214.480 380.280 215.600 ;
  LAYER ME2 ;
  RECT 376.740 214.480 380.280 215.600 ;
  LAYER ME1 ;
  RECT 376.740 214.480 380.280 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 368.060 214.480 371.600 215.600 ;
  LAYER ME3 ;
  RECT 368.060 214.480 371.600 215.600 ;
  LAYER ME2 ;
  RECT 368.060 214.480 371.600 215.600 ;
  LAYER ME1 ;
  RECT 368.060 214.480 371.600 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 359.380 214.480 362.920 215.600 ;
  LAYER ME3 ;
  RECT 359.380 214.480 362.920 215.600 ;
  LAYER ME2 ;
  RECT 359.380 214.480 362.920 215.600 ;
  LAYER ME1 ;
  RECT 359.380 214.480 362.920 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 315.980 214.480 319.520 215.600 ;
  LAYER ME3 ;
  RECT 315.980 214.480 319.520 215.600 ;
  LAYER ME2 ;
  RECT 315.980 214.480 319.520 215.600 ;
  LAYER ME1 ;
  RECT 315.980 214.480 319.520 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 307.300 214.480 310.840 215.600 ;
  LAYER ME3 ;
  RECT 307.300 214.480 310.840 215.600 ;
  LAYER ME2 ;
  RECT 307.300 214.480 310.840 215.600 ;
  LAYER ME1 ;
  RECT 307.300 214.480 310.840 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 298.620 214.480 302.160 215.600 ;
  LAYER ME3 ;
  RECT 298.620 214.480 302.160 215.600 ;
  LAYER ME2 ;
  RECT 298.620 214.480 302.160 215.600 ;
  LAYER ME1 ;
  RECT 298.620 214.480 302.160 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 289.940 214.480 293.480 215.600 ;
  LAYER ME3 ;
  RECT 289.940 214.480 293.480 215.600 ;
  LAYER ME2 ;
  RECT 289.940 214.480 293.480 215.600 ;
  LAYER ME1 ;
  RECT 289.940 214.480 293.480 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 281.260 214.480 284.800 215.600 ;
  LAYER ME3 ;
  RECT 281.260 214.480 284.800 215.600 ;
  LAYER ME2 ;
  RECT 281.260 214.480 284.800 215.600 ;
  LAYER ME1 ;
  RECT 281.260 214.480 284.800 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 272.580 214.480 276.120 215.600 ;
  LAYER ME3 ;
  RECT 272.580 214.480 276.120 215.600 ;
  LAYER ME2 ;
  RECT 272.580 214.480 276.120 215.600 ;
  LAYER ME1 ;
  RECT 272.580 214.480 276.120 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 229.180 214.480 232.720 215.600 ;
  LAYER ME3 ;
  RECT 229.180 214.480 232.720 215.600 ;
  LAYER ME2 ;
  RECT 229.180 214.480 232.720 215.600 ;
  LAYER ME1 ;
  RECT 229.180 214.480 232.720 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 220.500 214.480 224.040 215.600 ;
  LAYER ME3 ;
  RECT 220.500 214.480 224.040 215.600 ;
  LAYER ME2 ;
  RECT 220.500 214.480 224.040 215.600 ;
  LAYER ME1 ;
  RECT 220.500 214.480 224.040 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 211.820 214.480 215.360 215.600 ;
  LAYER ME3 ;
  RECT 211.820 214.480 215.360 215.600 ;
  LAYER ME2 ;
  RECT 211.820 214.480 215.360 215.600 ;
  LAYER ME1 ;
  RECT 211.820 214.480 215.360 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 203.140 214.480 206.680 215.600 ;
  LAYER ME3 ;
  RECT 203.140 214.480 206.680 215.600 ;
  LAYER ME2 ;
  RECT 203.140 214.480 206.680 215.600 ;
  LAYER ME1 ;
  RECT 203.140 214.480 206.680 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 194.460 214.480 198.000 215.600 ;
  LAYER ME3 ;
  RECT 194.460 214.480 198.000 215.600 ;
  LAYER ME2 ;
  RECT 194.460 214.480 198.000 215.600 ;
  LAYER ME1 ;
  RECT 194.460 214.480 198.000 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 185.780 214.480 189.320 215.600 ;
  LAYER ME3 ;
  RECT 185.780 214.480 189.320 215.600 ;
  LAYER ME2 ;
  RECT 185.780 214.480 189.320 215.600 ;
  LAYER ME1 ;
  RECT 185.780 214.480 189.320 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 142.380 214.480 145.920 215.600 ;
  LAYER ME3 ;
  RECT 142.380 214.480 145.920 215.600 ;
  LAYER ME2 ;
  RECT 142.380 214.480 145.920 215.600 ;
  LAYER ME1 ;
  RECT 142.380 214.480 145.920 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 133.700 214.480 137.240 215.600 ;
  LAYER ME3 ;
  RECT 133.700 214.480 137.240 215.600 ;
  LAYER ME2 ;
  RECT 133.700 214.480 137.240 215.600 ;
  LAYER ME1 ;
  RECT 133.700 214.480 137.240 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 125.020 214.480 128.560 215.600 ;
  LAYER ME3 ;
  RECT 125.020 214.480 128.560 215.600 ;
  LAYER ME2 ;
  RECT 125.020 214.480 128.560 215.600 ;
  LAYER ME1 ;
  RECT 125.020 214.480 128.560 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 116.340 214.480 119.880 215.600 ;
  LAYER ME3 ;
  RECT 116.340 214.480 119.880 215.600 ;
  LAYER ME2 ;
  RECT 116.340 214.480 119.880 215.600 ;
  LAYER ME1 ;
  RECT 116.340 214.480 119.880 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 107.660 214.480 111.200 215.600 ;
  LAYER ME3 ;
  RECT 107.660 214.480 111.200 215.600 ;
  LAYER ME2 ;
  RECT 107.660 214.480 111.200 215.600 ;
  LAYER ME1 ;
  RECT 107.660 214.480 111.200 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 98.980 214.480 102.520 215.600 ;
  LAYER ME3 ;
  RECT 98.980 214.480 102.520 215.600 ;
  LAYER ME2 ;
  RECT 98.980 214.480 102.520 215.600 ;
  LAYER ME1 ;
  RECT 98.980 214.480 102.520 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 55.580 214.480 59.120 215.600 ;
  LAYER ME3 ;
  RECT 55.580 214.480 59.120 215.600 ;
  LAYER ME2 ;
  RECT 55.580 214.480 59.120 215.600 ;
  LAYER ME1 ;
  RECT 55.580 214.480 59.120 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 46.900 214.480 50.440 215.600 ;
  LAYER ME3 ;
  RECT 46.900 214.480 50.440 215.600 ;
  LAYER ME2 ;
  RECT 46.900 214.480 50.440 215.600 ;
  LAYER ME1 ;
  RECT 46.900 214.480 50.440 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 38.220 214.480 41.760 215.600 ;
  LAYER ME3 ;
  RECT 38.220 214.480 41.760 215.600 ;
  LAYER ME2 ;
  RECT 38.220 214.480 41.760 215.600 ;
  LAYER ME1 ;
  RECT 38.220 214.480 41.760 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 29.540 214.480 33.080 215.600 ;
  LAYER ME3 ;
  RECT 29.540 214.480 33.080 215.600 ;
  LAYER ME2 ;
  RECT 29.540 214.480 33.080 215.600 ;
  LAYER ME1 ;
  RECT 29.540 214.480 33.080 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 20.860 214.480 24.400 215.600 ;
  LAYER ME3 ;
  RECT 20.860 214.480 24.400 215.600 ;
  LAYER ME2 ;
  RECT 20.860 214.480 24.400 215.600 ;
  LAYER ME1 ;
  RECT 20.860 214.480 24.400 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 12.180 214.480 15.720 215.600 ;
  LAYER ME3 ;
  RECT 12.180 214.480 15.720 215.600 ;
  LAYER ME2 ;
  RECT 12.180 214.480 15.720 215.600 ;
  LAYER ME1 ;
  RECT 12.180 214.480 15.720 215.600 ;
 END
 PORT
  LAYER ME4 ;
  RECT 531.120 0.000 534.660 1.120 ;
  LAYER ME3 ;
  RECT 531.120 0.000 534.660 1.120 ;
  LAYER ME2 ;
  RECT 531.120 0.000 534.660 1.120 ;
  LAYER ME1 ;
  RECT 531.120 0.000 534.660 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 509.420 0.000 512.960 1.120 ;
  LAYER ME3 ;
  RECT 509.420 0.000 512.960 1.120 ;
  LAYER ME2 ;
  RECT 509.420 0.000 512.960 1.120 ;
  LAYER ME1 ;
  RECT 509.420 0.000 512.960 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 492.680 0.000 496.220 1.120 ;
  LAYER ME3 ;
  RECT 492.680 0.000 496.220 1.120 ;
  LAYER ME2 ;
  RECT 492.680 0.000 496.220 1.120 ;
  LAYER ME1 ;
  RECT 492.680 0.000 496.220 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 466.020 0.000 469.560 1.120 ;
  LAYER ME3 ;
  RECT 466.020 0.000 469.560 1.120 ;
  LAYER ME2 ;
  RECT 466.020 0.000 469.560 1.120 ;
  LAYER ME1 ;
  RECT 466.020 0.000 469.560 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 353.180 0.000 356.720 1.120 ;
  LAYER ME3 ;
  RECT 353.180 0.000 356.720 1.120 ;
  LAYER ME2 ;
  RECT 353.180 0.000 356.720 1.120 ;
  LAYER ME1 ;
  RECT 353.180 0.000 356.720 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 331.480 0.000 335.020 1.120 ;
  LAYER ME3 ;
  RECT 331.480 0.000 335.020 1.120 ;
  LAYER ME2 ;
  RECT 331.480 0.000 335.020 1.120 ;
  LAYER ME1 ;
  RECT 331.480 0.000 335.020 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 309.780 0.000 313.320 1.120 ;
  LAYER ME3 ;
  RECT 309.780 0.000 313.320 1.120 ;
  LAYER ME2 ;
  RECT 309.780 0.000 313.320 1.120 ;
  LAYER ME1 ;
  RECT 309.780 0.000 313.320 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 282.500 0.000 286.040 1.120 ;
  LAYER ME3 ;
  RECT 282.500 0.000 286.040 1.120 ;
  LAYER ME2 ;
  RECT 282.500 0.000 286.040 1.120 ;
  LAYER ME1 ;
  RECT 282.500 0.000 286.040 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 273.820 0.000 277.360 1.120 ;
  LAYER ME3 ;
  RECT 273.820 0.000 277.360 1.120 ;
  LAYER ME2 ;
  RECT 273.820 0.000 277.360 1.120 ;
  LAYER ME1 ;
  RECT 273.820 0.000 277.360 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 246.540 0.000 250.080 1.120 ;
  LAYER ME3 ;
  RECT 246.540 0.000 250.080 1.120 ;
  LAYER ME2 ;
  RECT 246.540 0.000 250.080 1.120 ;
  LAYER ME1 ;
  RECT 246.540 0.000 250.080 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 139.900 0.000 143.440 1.120 ;
  LAYER ME3 ;
  RECT 139.900 0.000 143.440 1.120 ;
  LAYER ME2 ;
  RECT 139.900 0.000 143.440 1.120 ;
  LAYER ME1 ;
  RECT 139.900 0.000 143.440 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 113.860 0.000 117.400 1.120 ;
  LAYER ME3 ;
  RECT 113.860 0.000 117.400 1.120 ;
  LAYER ME2 ;
  RECT 113.860 0.000 117.400 1.120 ;
  LAYER ME1 ;
  RECT 113.860 0.000 117.400 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 92.160 0.000 95.700 1.120 ;
  LAYER ME3 ;
  RECT 92.160 0.000 95.700 1.120 ;
  LAYER ME2 ;
  RECT 92.160 0.000 95.700 1.120 ;
  LAYER ME1 ;
  RECT 92.160 0.000 95.700 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 70.460 0.000 74.000 1.120 ;
  LAYER ME3 ;
  RECT 70.460 0.000 74.000 1.120 ;
  LAYER ME2 ;
  RECT 70.460 0.000 74.000 1.120 ;
  LAYER ME1 ;
  RECT 70.460 0.000 74.000 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 43.800 0.000 47.340 1.120 ;
  LAYER ME3 ;
  RECT 43.800 0.000 47.340 1.120 ;
  LAYER ME2 ;
  RECT 43.800 0.000 47.340 1.120 ;
  LAYER ME1 ;
  RECT 43.800 0.000 47.340 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 27.060 0.000 30.600 1.120 ;
  LAYER ME3 ;
  RECT 27.060 0.000 30.600 1.120 ;
  LAYER ME2 ;
  RECT 27.060 0.000 30.600 1.120 ;
  LAYER ME1 ;
  RECT 27.060 0.000 30.600 1.120 ;
 END
END GND
PIN DO31
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 528.920 0.000 530.040 1.120 ;
  LAYER ME3 ;
  RECT 528.920 0.000 530.040 1.120 ;
  LAYER ME2 ;
  RECT 528.920 0.000 530.040 1.120 ;
  LAYER ME1 ;
  RECT 528.920 0.000 530.040 1.120 ;
 END
END DO31
PIN DI31
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 520.240 0.000 521.360 1.120 ;
  LAYER ME3 ;
  RECT 520.240 0.000 521.360 1.120 ;
  LAYER ME2 ;
  RECT 520.240 0.000 521.360 1.120 ;
  LAYER ME1 ;
  RECT 520.240 0.000 521.360 1.120 ;
 END
END DI31
PIN DO30
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 515.280 0.000 516.400 1.120 ;
  LAYER ME3 ;
  RECT 515.280 0.000 516.400 1.120 ;
  LAYER ME2 ;
  RECT 515.280 0.000 516.400 1.120 ;
  LAYER ME1 ;
  RECT 515.280 0.000 516.400 1.120 ;
 END
END DO30
PIN DI30
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 507.220 0.000 508.340 1.120 ;
  LAYER ME3 ;
  RECT 507.220 0.000 508.340 1.120 ;
  LAYER ME2 ;
  RECT 507.220 0.000 508.340 1.120 ;
  LAYER ME1 ;
  RECT 507.220 0.000 508.340 1.120 ;
 END
END DI30
PIN DO29
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 498.540 0.000 499.660 1.120 ;
  LAYER ME3 ;
  RECT 498.540 0.000 499.660 1.120 ;
  LAYER ME2 ;
  RECT 498.540 0.000 499.660 1.120 ;
  LAYER ME1 ;
  RECT 498.540 0.000 499.660 1.120 ;
 END
END DO29
PIN DI29
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 490.480 0.000 491.600 1.120 ;
  LAYER ME3 ;
  RECT 490.480 0.000 491.600 1.120 ;
  LAYER ME2 ;
  RECT 490.480 0.000 491.600 1.120 ;
  LAYER ME1 ;
  RECT 490.480 0.000 491.600 1.120 ;
 END
END DI29
PIN DO28
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 485.520 0.000 486.640 1.120 ;
  LAYER ME3 ;
  RECT 485.520 0.000 486.640 1.120 ;
  LAYER ME2 ;
  RECT 485.520 0.000 486.640 1.120 ;
  LAYER ME1 ;
  RECT 485.520 0.000 486.640 1.120 ;
 END
END DO28
PIN DI28
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 477.460 0.000 478.580 1.120 ;
  LAYER ME3 ;
  RECT 477.460 0.000 478.580 1.120 ;
  LAYER ME2 ;
  RECT 477.460 0.000 478.580 1.120 ;
  LAYER ME1 ;
  RECT 477.460 0.000 478.580 1.120 ;
 END
END DI28
PIN DO27
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 472.500 0.000 473.620 1.120 ;
  LAYER ME3 ;
  RECT 472.500 0.000 473.620 1.120 ;
  LAYER ME2 ;
  RECT 472.500 0.000 473.620 1.120 ;
  LAYER ME1 ;
  RECT 472.500 0.000 473.620 1.120 ;
 END
END DO27
PIN DI27
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 463.820 0.000 464.940 1.120 ;
  LAYER ME3 ;
  RECT 463.820 0.000 464.940 1.120 ;
  LAYER ME2 ;
  RECT 463.820 0.000 464.940 1.120 ;
  LAYER ME1 ;
  RECT 463.820 0.000 464.940 1.120 ;
 END
END DI27
PIN DO26
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 458.860 0.000 459.980 1.120 ;
  LAYER ME3 ;
  RECT 458.860 0.000 459.980 1.120 ;
  LAYER ME2 ;
  RECT 458.860 0.000 459.980 1.120 ;
  LAYER ME1 ;
  RECT 458.860 0.000 459.980 1.120 ;
 END
END DO26
PIN DI26
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 450.800 0.000 451.920 1.120 ;
  LAYER ME3 ;
  RECT 450.800 0.000 451.920 1.120 ;
  LAYER ME2 ;
  RECT 450.800 0.000 451.920 1.120 ;
  LAYER ME1 ;
  RECT 450.800 0.000 451.920 1.120 ;
 END
END DI26
PIN DO25
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 442.120 0.000 443.240 1.120 ;
  LAYER ME3 ;
  RECT 442.120 0.000 443.240 1.120 ;
  LAYER ME2 ;
  RECT 442.120 0.000 443.240 1.120 ;
  LAYER ME1 ;
  RECT 442.120 0.000 443.240 1.120 ;
 END
END DO25
PIN DI25
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 434.060 0.000 435.180 1.120 ;
  LAYER ME3 ;
  RECT 434.060 0.000 435.180 1.120 ;
  LAYER ME2 ;
  RECT 434.060 0.000 435.180 1.120 ;
  LAYER ME1 ;
  RECT 434.060 0.000 435.180 1.120 ;
 END
END DI25
PIN DO24
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 429.100 0.000 430.220 1.120 ;
  LAYER ME3 ;
  RECT 429.100 0.000 430.220 1.120 ;
  LAYER ME2 ;
  RECT 429.100 0.000 430.220 1.120 ;
  LAYER ME1 ;
  RECT 429.100 0.000 430.220 1.120 ;
 END
END DO24
PIN DI24
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 420.420 0.000 421.540 1.120 ;
  LAYER ME3 ;
  RECT 420.420 0.000 421.540 1.120 ;
  LAYER ME2 ;
  RECT 420.420 0.000 421.540 1.120 ;
  LAYER ME1 ;
  RECT 420.420 0.000 421.540 1.120 ;
 END
END DI24
PIN DO23
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 415.460 0.000 416.580 1.120 ;
  LAYER ME3 ;
  RECT 415.460 0.000 416.580 1.120 ;
  LAYER ME2 ;
  RECT 415.460 0.000 416.580 1.120 ;
  LAYER ME1 ;
  RECT 415.460 0.000 416.580 1.120 ;
 END
END DO23
PIN DI23
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 407.400 0.000 408.520 1.120 ;
  LAYER ME3 ;
  RECT 407.400 0.000 408.520 1.120 ;
  LAYER ME2 ;
  RECT 407.400 0.000 408.520 1.120 ;
  LAYER ME1 ;
  RECT 407.400 0.000 408.520 1.120 ;
 END
END DI23
PIN DO22
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 402.440 0.000 403.560 1.120 ;
  LAYER ME3 ;
  RECT 402.440 0.000 403.560 1.120 ;
  LAYER ME2 ;
  RECT 402.440 0.000 403.560 1.120 ;
  LAYER ME1 ;
  RECT 402.440 0.000 403.560 1.120 ;
 END
END DO22
PIN DI22
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 394.380 0.000 395.500 1.120 ;
  LAYER ME3 ;
  RECT 394.380 0.000 395.500 1.120 ;
  LAYER ME2 ;
  RECT 394.380 0.000 395.500 1.120 ;
  LAYER ME1 ;
  RECT 394.380 0.000 395.500 1.120 ;
 END
END DI22
PIN DO21
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 385.700 0.000 386.820 1.120 ;
  LAYER ME3 ;
  RECT 385.700 0.000 386.820 1.120 ;
  LAYER ME2 ;
  RECT 385.700 0.000 386.820 1.120 ;
  LAYER ME1 ;
  RECT 385.700 0.000 386.820 1.120 ;
 END
END DO21
PIN DI21
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 377.640 0.000 378.760 1.120 ;
  LAYER ME3 ;
  RECT 377.640 0.000 378.760 1.120 ;
  LAYER ME2 ;
  RECT 377.640 0.000 378.760 1.120 ;
  LAYER ME1 ;
  RECT 377.640 0.000 378.760 1.120 ;
 END
END DI21
PIN DO20
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 372.680 0.000 373.800 1.120 ;
  LAYER ME3 ;
  RECT 372.680 0.000 373.800 1.120 ;
  LAYER ME2 ;
  RECT 372.680 0.000 373.800 1.120 ;
  LAYER ME1 ;
  RECT 372.680 0.000 373.800 1.120 ;
 END
END DO20
PIN DI20
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 364.000 0.000 365.120 1.120 ;
  LAYER ME3 ;
  RECT 364.000 0.000 365.120 1.120 ;
  LAYER ME2 ;
  RECT 364.000 0.000 365.120 1.120 ;
  LAYER ME1 ;
  RECT 364.000 0.000 365.120 1.120 ;
 END
END DI20
PIN DO19
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 359.040 0.000 360.160 1.120 ;
  LAYER ME3 ;
  RECT 359.040 0.000 360.160 1.120 ;
  LAYER ME2 ;
  RECT 359.040 0.000 360.160 1.120 ;
  LAYER ME1 ;
  RECT 359.040 0.000 360.160 1.120 ;
 END
END DO19
PIN DI19
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 350.980 0.000 352.100 1.120 ;
  LAYER ME3 ;
  RECT 350.980 0.000 352.100 1.120 ;
  LAYER ME2 ;
  RECT 350.980 0.000 352.100 1.120 ;
  LAYER ME1 ;
  RECT 350.980 0.000 352.100 1.120 ;
 END
END DI19
PIN DO18
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 346.020 0.000 347.140 1.120 ;
  LAYER ME3 ;
  RECT 346.020 0.000 347.140 1.120 ;
  LAYER ME2 ;
  RECT 346.020 0.000 347.140 1.120 ;
  LAYER ME1 ;
  RECT 346.020 0.000 347.140 1.120 ;
 END
END DO18
PIN DI18
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 337.340 0.000 338.460 1.120 ;
  LAYER ME3 ;
  RECT 337.340 0.000 338.460 1.120 ;
  LAYER ME2 ;
  RECT 337.340 0.000 338.460 1.120 ;
  LAYER ME1 ;
  RECT 337.340 0.000 338.460 1.120 ;
 END
END DI18
PIN DO17
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 329.280 0.000 330.400 1.120 ;
  LAYER ME3 ;
  RECT 329.280 0.000 330.400 1.120 ;
  LAYER ME2 ;
  RECT 329.280 0.000 330.400 1.120 ;
  LAYER ME1 ;
  RECT 329.280 0.000 330.400 1.120 ;
 END
END DO17
PIN DI17
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 320.600 0.000 321.720 1.120 ;
  LAYER ME3 ;
  RECT 320.600 0.000 321.720 1.120 ;
  LAYER ME2 ;
  RECT 320.600 0.000 321.720 1.120 ;
  LAYER ME1 ;
  RECT 320.600 0.000 321.720 1.120 ;
 END
END DI17
PIN DO16
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 316.260 0.000 317.380 1.120 ;
  LAYER ME3 ;
  RECT 316.260 0.000 317.380 1.120 ;
  LAYER ME2 ;
  RECT 316.260 0.000 317.380 1.120 ;
  LAYER ME1 ;
  RECT 316.260 0.000 317.380 1.120 ;
 END
END DO16
PIN DI16
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 307.580 0.000 308.700 1.120 ;
  LAYER ME3 ;
  RECT 307.580 0.000 308.700 1.120 ;
  LAYER ME2 ;
  RECT 307.580 0.000 308.700 1.120 ;
  LAYER ME1 ;
  RECT 307.580 0.000 308.700 1.120 ;
 END
END DI16
PIN A1
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 302.000 0.000 303.120 1.120 ;
  LAYER ME3 ;
  RECT 302.000 0.000 303.120 1.120 ;
  LAYER ME2 ;
  RECT 302.000 0.000 303.120 1.120 ;
  LAYER ME1 ;
  RECT 302.000 0.000 303.120 1.120 ;
 END
END A1
PIN WEB
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER ME4 ;
  RECT 300.140 0.000 301.260 1.120 ;
  LAYER ME3 ;
  RECT 300.140 0.000 301.260 1.120 ;
  LAYER ME2 ;
  RECT 300.140 0.000 301.260 1.120 ;
  LAYER ME1 ;
  RECT 300.140 0.000 301.260 1.120 ;
 END
END WEB
PIN OE
  DIRECTION INPUT ;
  CAPACITANCE 0.033 ;
 PORT
  LAYER ME4 ;
  RECT 295.180 0.000 296.300 1.120 ;
  LAYER ME3 ;
  RECT 295.180 0.000 296.300 1.120 ;
  LAYER ME2 ;
  RECT 295.180 0.000 296.300 1.120 ;
  LAYER ME1 ;
  RECT 295.180 0.000 296.300 1.120 ;
 END
END OE
PIN CS
  DIRECTION INPUT ;
  CAPACITANCE 0.123 ;
 PORT
  LAYER ME4 ;
  RECT 293.320 0.000 294.440 1.120 ;
  LAYER ME3 ;
  RECT 293.320 0.000 294.440 1.120 ;
  LAYER ME2 ;
  RECT 293.320 0.000 294.440 1.120 ;
  LAYER ME1 ;
  RECT 293.320 0.000 294.440 1.120 ;
 END
END CS
PIN A2
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 271.620 0.000 272.740 1.120 ;
  LAYER ME3 ;
  RECT 271.620 0.000 272.740 1.120 ;
  LAYER ME2 ;
  RECT 271.620 0.000 272.740 1.120 ;
  LAYER ME1 ;
  RECT 271.620 0.000 272.740 1.120 ;
 END
END A2
PIN CK
  DIRECTION INPUT ;
  CAPACITANCE 0.063 ;
 PORT
  LAYER ME4 ;
  RECT 268.520 0.000 269.640 1.120 ;
  LAYER ME3 ;
  RECT 268.520 0.000 269.640 1.120 ;
  LAYER ME2 ;
  RECT 268.520 0.000 269.640 1.120 ;
  LAYER ME1 ;
  RECT 268.520 0.000 269.640 1.120 ;
 END
END CK
PIN A0
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 266.660 0.000 267.780 1.120 ;
  LAYER ME3 ;
  RECT 266.660 0.000 267.780 1.120 ;
  LAYER ME2 ;
  RECT 266.660 0.000 267.780 1.120 ;
  LAYER ME1 ;
  RECT 266.660 0.000 267.780 1.120 ;
 END
END A0
PIN A3
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 262.320 0.000 263.440 1.120 ;
  LAYER ME3 ;
  RECT 262.320 0.000 263.440 1.120 ;
  LAYER ME2 ;
  RECT 262.320 0.000 263.440 1.120 ;
  LAYER ME1 ;
  RECT 262.320 0.000 263.440 1.120 ;
 END
END A3
PIN A4
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 254.880 0.000 256.000 1.120 ;
  LAYER ME3 ;
  RECT 254.880 0.000 256.000 1.120 ;
  LAYER ME2 ;
  RECT 254.880 0.000 256.000 1.120 ;
  LAYER ME1 ;
  RECT 254.880 0.000 256.000 1.120 ;
 END
END A4
PIN A5
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 251.780 0.000 252.900 1.120 ;
  LAYER ME3 ;
  RECT 251.780 0.000 252.900 1.120 ;
  LAYER ME2 ;
  RECT 251.780 0.000 252.900 1.120 ;
  LAYER ME1 ;
  RECT 251.780 0.000 252.900 1.120 ;
 END
END A5
PIN A6
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 244.340 0.000 245.460 1.120 ;
  LAYER ME3 ;
  RECT 244.340 0.000 245.460 1.120 ;
  LAYER ME2 ;
  RECT 244.340 0.000 245.460 1.120 ;
  LAYER ME1 ;
  RECT 244.340 0.000 245.460 1.120 ;
 END
END A6
PIN A7
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 241.240 0.000 242.360 1.120 ;
  LAYER ME3 ;
  RECT 241.240 0.000 242.360 1.120 ;
  LAYER ME2 ;
  RECT 241.240 0.000 242.360 1.120 ;
  LAYER ME1 ;
  RECT 241.240 0.000 242.360 1.120 ;
 END
END A7
PIN DO15
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 233.180 0.000 234.300 1.120 ;
  LAYER ME3 ;
  RECT 233.180 0.000 234.300 1.120 ;
  LAYER ME2 ;
  RECT 233.180 0.000 234.300 1.120 ;
  LAYER ME1 ;
  RECT 233.180 0.000 234.300 1.120 ;
 END
END DO15
PIN DI15
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 224.500 0.000 225.620 1.120 ;
  LAYER ME3 ;
  RECT 224.500 0.000 225.620 1.120 ;
  LAYER ME2 ;
  RECT 224.500 0.000 225.620 1.120 ;
  LAYER ME1 ;
  RECT 224.500 0.000 225.620 1.120 ;
 END
END DI15
PIN DO14
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 219.540 0.000 220.660 1.120 ;
  LAYER ME3 ;
  RECT 219.540 0.000 220.660 1.120 ;
  LAYER ME2 ;
  RECT 219.540 0.000 220.660 1.120 ;
  LAYER ME1 ;
  RECT 219.540 0.000 220.660 1.120 ;
 END
END DO14
PIN DI14
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 211.480 0.000 212.600 1.120 ;
  LAYER ME3 ;
  RECT 211.480 0.000 212.600 1.120 ;
  LAYER ME2 ;
  RECT 211.480 0.000 212.600 1.120 ;
  LAYER ME1 ;
  RECT 211.480 0.000 212.600 1.120 ;
 END
END DI14
PIN DO13
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 202.800 0.000 203.920 1.120 ;
  LAYER ME3 ;
  RECT 202.800 0.000 203.920 1.120 ;
  LAYER ME2 ;
  RECT 202.800 0.000 203.920 1.120 ;
  LAYER ME1 ;
  RECT 202.800 0.000 203.920 1.120 ;
 END
END DO13
PIN DI13
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 194.740 0.000 195.860 1.120 ;
  LAYER ME3 ;
  RECT 194.740 0.000 195.860 1.120 ;
  LAYER ME2 ;
  RECT 194.740 0.000 195.860 1.120 ;
  LAYER ME1 ;
  RECT 194.740 0.000 195.860 1.120 ;
 END
END DI13
PIN DO12
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 189.780 0.000 190.900 1.120 ;
  LAYER ME3 ;
  RECT 189.780 0.000 190.900 1.120 ;
  LAYER ME2 ;
  RECT 189.780 0.000 190.900 1.120 ;
  LAYER ME1 ;
  RECT 189.780 0.000 190.900 1.120 ;
 END
END DO12
PIN DI12
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 181.100 0.000 182.220 1.120 ;
  LAYER ME3 ;
  RECT 181.100 0.000 182.220 1.120 ;
  LAYER ME2 ;
  RECT 181.100 0.000 182.220 1.120 ;
  LAYER ME1 ;
  RECT 181.100 0.000 182.220 1.120 ;
 END
END DI12
PIN DO11
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 176.140 0.000 177.260 1.120 ;
  LAYER ME3 ;
  RECT 176.140 0.000 177.260 1.120 ;
  LAYER ME2 ;
  RECT 176.140 0.000 177.260 1.120 ;
  LAYER ME1 ;
  RECT 176.140 0.000 177.260 1.120 ;
 END
END DO11
PIN DI11
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 168.080 0.000 169.200 1.120 ;
  LAYER ME3 ;
  RECT 168.080 0.000 169.200 1.120 ;
  LAYER ME2 ;
  RECT 168.080 0.000 169.200 1.120 ;
  LAYER ME1 ;
  RECT 168.080 0.000 169.200 1.120 ;
 END
END DI11
PIN DO10
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 163.120 0.000 164.240 1.120 ;
  LAYER ME3 ;
  RECT 163.120 0.000 164.240 1.120 ;
  LAYER ME2 ;
  RECT 163.120 0.000 164.240 1.120 ;
  LAYER ME1 ;
  RECT 163.120 0.000 164.240 1.120 ;
 END
END DO10
PIN DI10
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 154.440 0.000 155.560 1.120 ;
  LAYER ME3 ;
  RECT 154.440 0.000 155.560 1.120 ;
  LAYER ME2 ;
  RECT 154.440 0.000 155.560 1.120 ;
  LAYER ME1 ;
  RECT 154.440 0.000 155.560 1.120 ;
 END
END DI10
PIN DO9
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 146.380 0.000 147.500 1.120 ;
  LAYER ME3 ;
  RECT 146.380 0.000 147.500 1.120 ;
  LAYER ME2 ;
  RECT 146.380 0.000 147.500 1.120 ;
  LAYER ME1 ;
  RECT 146.380 0.000 147.500 1.120 ;
 END
END DO9
PIN DI9
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 137.700 0.000 138.820 1.120 ;
  LAYER ME3 ;
  RECT 137.700 0.000 138.820 1.120 ;
  LAYER ME2 ;
  RECT 137.700 0.000 138.820 1.120 ;
  LAYER ME1 ;
  RECT 137.700 0.000 138.820 1.120 ;
 END
END DI9
PIN DO8
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 133.360 0.000 134.480 1.120 ;
  LAYER ME3 ;
  RECT 133.360 0.000 134.480 1.120 ;
  LAYER ME2 ;
  RECT 133.360 0.000 134.480 1.120 ;
  LAYER ME1 ;
  RECT 133.360 0.000 134.480 1.120 ;
 END
END DO8
PIN DI8
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 124.680 0.000 125.800 1.120 ;
  LAYER ME3 ;
  RECT 124.680 0.000 125.800 1.120 ;
  LAYER ME2 ;
  RECT 124.680 0.000 125.800 1.120 ;
  LAYER ME1 ;
  RECT 124.680 0.000 125.800 1.120 ;
 END
END DI8
PIN DO7
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 119.720 0.000 120.840 1.120 ;
  LAYER ME3 ;
  RECT 119.720 0.000 120.840 1.120 ;
  LAYER ME2 ;
  RECT 119.720 0.000 120.840 1.120 ;
  LAYER ME1 ;
  RECT 119.720 0.000 120.840 1.120 ;
 END
END DO7
PIN DI7
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 111.660 0.000 112.780 1.120 ;
  LAYER ME3 ;
  RECT 111.660 0.000 112.780 1.120 ;
  LAYER ME2 ;
  RECT 111.660 0.000 112.780 1.120 ;
  LAYER ME1 ;
  RECT 111.660 0.000 112.780 1.120 ;
 END
END DI7
PIN DO6
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 106.700 0.000 107.820 1.120 ;
  LAYER ME3 ;
  RECT 106.700 0.000 107.820 1.120 ;
  LAYER ME2 ;
  RECT 106.700 0.000 107.820 1.120 ;
  LAYER ME1 ;
  RECT 106.700 0.000 107.820 1.120 ;
 END
END DO6
PIN DI6
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 98.020 0.000 99.140 1.120 ;
  LAYER ME3 ;
  RECT 98.020 0.000 99.140 1.120 ;
  LAYER ME2 ;
  RECT 98.020 0.000 99.140 1.120 ;
  LAYER ME1 ;
  RECT 98.020 0.000 99.140 1.120 ;
 END
END DI6
PIN DO5
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 89.960 0.000 91.080 1.120 ;
  LAYER ME3 ;
  RECT 89.960 0.000 91.080 1.120 ;
  LAYER ME2 ;
  RECT 89.960 0.000 91.080 1.120 ;
  LAYER ME1 ;
  RECT 89.960 0.000 91.080 1.120 ;
 END
END DO5
PIN DI5
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 81.280 0.000 82.400 1.120 ;
  LAYER ME3 ;
  RECT 81.280 0.000 82.400 1.120 ;
  LAYER ME2 ;
  RECT 81.280 0.000 82.400 1.120 ;
  LAYER ME1 ;
  RECT 81.280 0.000 82.400 1.120 ;
 END
END DI5
PIN DO4
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 76.320 0.000 77.440 1.120 ;
  LAYER ME3 ;
  RECT 76.320 0.000 77.440 1.120 ;
  LAYER ME2 ;
  RECT 76.320 0.000 77.440 1.120 ;
  LAYER ME1 ;
  RECT 76.320 0.000 77.440 1.120 ;
 END
END DO4
PIN DI4
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 68.260 0.000 69.380 1.120 ;
  LAYER ME3 ;
  RECT 68.260 0.000 69.380 1.120 ;
  LAYER ME2 ;
  RECT 68.260 0.000 69.380 1.120 ;
  LAYER ME1 ;
  RECT 68.260 0.000 69.380 1.120 ;
 END
END DI4
PIN DO3
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 63.300 0.000 64.420 1.120 ;
  LAYER ME3 ;
  RECT 63.300 0.000 64.420 1.120 ;
  LAYER ME2 ;
  RECT 63.300 0.000 64.420 1.120 ;
  LAYER ME1 ;
  RECT 63.300 0.000 64.420 1.120 ;
 END
END DO3
PIN DI3
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 54.620 0.000 55.740 1.120 ;
  LAYER ME3 ;
  RECT 54.620 0.000 55.740 1.120 ;
  LAYER ME2 ;
  RECT 54.620 0.000 55.740 1.120 ;
  LAYER ME1 ;
  RECT 54.620 0.000 55.740 1.120 ;
 END
END DI3
PIN DO2
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 50.280 0.000 51.400 1.120 ;
  LAYER ME3 ;
  RECT 50.280 0.000 51.400 1.120 ;
  LAYER ME2 ;
  RECT 50.280 0.000 51.400 1.120 ;
  LAYER ME1 ;
  RECT 50.280 0.000 51.400 1.120 ;
 END
END DO2
PIN DI2
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 41.600 0.000 42.720 1.120 ;
  LAYER ME3 ;
  RECT 41.600 0.000 42.720 1.120 ;
  LAYER ME2 ;
  RECT 41.600 0.000 42.720 1.120 ;
  LAYER ME1 ;
  RECT 41.600 0.000 42.720 1.120 ;
 END
END DI2
PIN DO1
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 33.540 0.000 34.660 1.120 ;
  LAYER ME3 ;
  RECT 33.540 0.000 34.660 1.120 ;
  LAYER ME2 ;
  RECT 33.540 0.000 34.660 1.120 ;
  LAYER ME1 ;
  RECT 33.540 0.000 34.660 1.120 ;
 END
END DO1
PIN DI1
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 24.860 0.000 25.980 1.120 ;
  LAYER ME3 ;
  RECT 24.860 0.000 25.980 1.120 ;
  LAYER ME2 ;
  RECT 24.860 0.000 25.980 1.120 ;
  LAYER ME1 ;
  RECT 24.860 0.000 25.980 1.120 ;
 END
END DI1
PIN DO0
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 19.900 0.000 21.020 1.120 ;
  LAYER ME3 ;
  RECT 19.900 0.000 21.020 1.120 ;
  LAYER ME2 ;
  RECT 19.900 0.000 21.020 1.120 ;
  LAYER ME1 ;
  RECT 19.900 0.000 21.020 1.120 ;
 END
END DO0
PIN DI0
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 11.840 0.000 12.960 1.120 ;
  LAYER ME3 ;
  RECT 11.840 0.000 12.960 1.120 ;
  LAYER ME2 ;
  RECT 11.840 0.000 12.960 1.120 ;
  LAYER ME1 ;
  RECT 11.840 0.000 12.960 1.120 ;
 END
END DI0
OBS
  LAYER ME1 SPACING 0.280 ;
  RECT 0.000 0.140 542.500 215.600 ;
  LAYER ME2 SPACING 0.320 ;
  RECT 0.000 0.140 542.500 215.600 ;
  LAYER ME3 SPACING 0.320 ;
  RECT 0.000 0.140 542.500 215.600 ;
  LAYER ME4 SPACING 0.600 ;
  RECT 0.000 0.140 542.500 215.600 ;
  LAYER VI1 ;
  RECT 0.000 0.140 542.500 215.600 ;
  LAYER VI2 ;
  RECT 0.000 0.140 542.500 215.600 ;
  LAYER VI3 ;
  RECT 0.000 0.140 542.500 215.600 ;
END
END Memory_32_256
END LIBRARY



