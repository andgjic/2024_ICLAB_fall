# 
#              Synchronous High Speed Single Port SRAM Compiler 
# 
#                    UMC 0.18um GenericII Logic Process
#    __________________________________________________________________________
# 
# 
#      (C) Copyright 2002-2009 Faraday Technology Corp. All Rights Reserved.
#    
#    This source code is an unpublished work belongs to Faraday Technology
#    Corp.  It is considered a trade secret and is not to be divulged or
#    used by parties who have not received written authorization from
#    Faraday Technology Corp.
#    
#    Faraday's home page can be found at:
#    http://www.faraday-tech.com/
#   
#       Module Name      : Memory_64_128
#       Words            : 128
#       Bits             : 64
#       Byte-Write       : 1
#       Aspect Ratio     : 1
#       Output Loading   : 0.05  (pf)
#       Data Slew        : 0.02  (ns)
#       CK Slew          : 0.02  (ns)
#       Power Ring Width : 2  (um)
# 
# -----------------------------------------------------------------------------
# 
#       Library          : FSA0M_A
#       Memaker          : 200901.2.1
#       Date             : 2024/10/27 11:40:58
# 
# -----------------------------------------------------------------------------


NAMESCASESENSITIVE ON ;
MACRO Memory_64_128
CLASS BLOCK ;
FOREIGN Memory_64_128 0.000 0.000 ;
ORIGIN 0.000 0.000 ;
SIZE 994.480 BY 176.400 ;
SYMMETRY x y r90 ;
SITE core ;
PIN VCC
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
 PORT
  LAYER ME4 ;
  RECT 993.360 164.980 994.480 168.220 ;
  LAYER ME3 ;
  RECT 993.360 164.980 994.480 168.220 ;
  LAYER ME2 ;
  RECT 993.360 164.980 994.480 168.220 ;
  LAYER ME1 ;
  RECT 993.360 164.980 994.480 168.220 ;
 END
 PORT
  LAYER ME4 ;
  RECT 993.360 125.780 994.480 129.020 ;
  LAYER ME3 ;
  RECT 993.360 125.780 994.480 129.020 ;
  LAYER ME2 ;
  RECT 993.360 125.780 994.480 129.020 ;
  LAYER ME1 ;
  RECT 993.360 125.780 994.480 129.020 ;
 END
 PORT
  LAYER ME4 ;
  RECT 993.360 117.940 994.480 121.180 ;
  LAYER ME3 ;
  RECT 993.360 117.940 994.480 121.180 ;
  LAYER ME2 ;
  RECT 993.360 117.940 994.480 121.180 ;
  LAYER ME1 ;
  RECT 993.360 117.940 994.480 121.180 ;
 END
 PORT
  LAYER ME4 ;
  RECT 993.360 110.100 994.480 113.340 ;
  LAYER ME3 ;
  RECT 993.360 110.100 994.480 113.340 ;
  LAYER ME2 ;
  RECT 993.360 110.100 994.480 113.340 ;
  LAYER ME1 ;
  RECT 993.360 110.100 994.480 113.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 993.360 102.260 994.480 105.500 ;
  LAYER ME3 ;
  RECT 993.360 102.260 994.480 105.500 ;
  LAYER ME2 ;
  RECT 993.360 102.260 994.480 105.500 ;
  LAYER ME1 ;
  RECT 993.360 102.260 994.480 105.500 ;
 END
 PORT
  LAYER ME4 ;
  RECT 993.360 94.420 994.480 97.660 ;
  LAYER ME3 ;
  RECT 993.360 94.420 994.480 97.660 ;
  LAYER ME2 ;
  RECT 993.360 94.420 994.480 97.660 ;
  LAYER ME1 ;
  RECT 993.360 94.420 994.480 97.660 ;
 END
 PORT
  LAYER ME4 ;
  RECT 993.360 86.580 994.480 89.820 ;
  LAYER ME3 ;
  RECT 993.360 86.580 994.480 89.820 ;
  LAYER ME2 ;
  RECT 993.360 86.580 994.480 89.820 ;
  LAYER ME1 ;
  RECT 993.360 86.580 994.480 89.820 ;
 END
 PORT
  LAYER ME4 ;
  RECT 993.360 47.380 994.480 50.620 ;
  LAYER ME3 ;
  RECT 993.360 47.380 994.480 50.620 ;
  LAYER ME2 ;
  RECT 993.360 47.380 994.480 50.620 ;
  LAYER ME1 ;
  RECT 993.360 47.380 994.480 50.620 ;
 END
 PORT
  LAYER ME4 ;
  RECT 993.360 39.540 994.480 42.780 ;
  LAYER ME3 ;
  RECT 993.360 39.540 994.480 42.780 ;
  LAYER ME2 ;
  RECT 993.360 39.540 994.480 42.780 ;
  LAYER ME1 ;
  RECT 993.360 39.540 994.480 42.780 ;
 END
 PORT
  LAYER ME4 ;
  RECT 993.360 31.700 994.480 34.940 ;
  LAYER ME3 ;
  RECT 993.360 31.700 994.480 34.940 ;
  LAYER ME2 ;
  RECT 993.360 31.700 994.480 34.940 ;
  LAYER ME1 ;
  RECT 993.360 31.700 994.480 34.940 ;
 END
 PORT
  LAYER ME4 ;
  RECT 993.360 23.860 994.480 27.100 ;
  LAYER ME3 ;
  RECT 993.360 23.860 994.480 27.100 ;
  LAYER ME2 ;
  RECT 993.360 23.860 994.480 27.100 ;
  LAYER ME1 ;
  RECT 993.360 23.860 994.480 27.100 ;
 END
 PORT
  LAYER ME4 ;
  RECT 993.360 16.020 994.480 19.260 ;
  LAYER ME3 ;
  RECT 993.360 16.020 994.480 19.260 ;
  LAYER ME2 ;
  RECT 993.360 16.020 994.480 19.260 ;
  LAYER ME1 ;
  RECT 993.360 16.020 994.480 19.260 ;
 END
 PORT
  LAYER ME4 ;
  RECT 993.360 8.180 994.480 11.420 ;
  LAYER ME3 ;
  RECT 993.360 8.180 994.480 11.420 ;
  LAYER ME2 ;
  RECT 993.360 8.180 994.480 11.420 ;
  LAYER ME1 ;
  RECT 993.360 8.180 994.480 11.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 164.980 1.120 168.220 ;
  LAYER ME3 ;
  RECT 0.000 164.980 1.120 168.220 ;
  LAYER ME2 ;
  RECT 0.000 164.980 1.120 168.220 ;
  LAYER ME1 ;
  RECT 0.000 164.980 1.120 168.220 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 125.780 1.120 129.020 ;
  LAYER ME3 ;
  RECT 0.000 125.780 1.120 129.020 ;
  LAYER ME2 ;
  RECT 0.000 125.780 1.120 129.020 ;
  LAYER ME1 ;
  RECT 0.000 125.780 1.120 129.020 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 117.940 1.120 121.180 ;
  LAYER ME3 ;
  RECT 0.000 117.940 1.120 121.180 ;
  LAYER ME2 ;
  RECT 0.000 117.940 1.120 121.180 ;
  LAYER ME1 ;
  RECT 0.000 117.940 1.120 121.180 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 110.100 1.120 113.340 ;
  LAYER ME3 ;
  RECT 0.000 110.100 1.120 113.340 ;
  LAYER ME2 ;
  RECT 0.000 110.100 1.120 113.340 ;
  LAYER ME1 ;
  RECT 0.000 110.100 1.120 113.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 102.260 1.120 105.500 ;
  LAYER ME3 ;
  RECT 0.000 102.260 1.120 105.500 ;
  LAYER ME2 ;
  RECT 0.000 102.260 1.120 105.500 ;
  LAYER ME1 ;
  RECT 0.000 102.260 1.120 105.500 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 94.420 1.120 97.660 ;
  LAYER ME3 ;
  RECT 0.000 94.420 1.120 97.660 ;
  LAYER ME2 ;
  RECT 0.000 94.420 1.120 97.660 ;
  LAYER ME1 ;
  RECT 0.000 94.420 1.120 97.660 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 86.580 1.120 89.820 ;
  LAYER ME3 ;
  RECT 0.000 86.580 1.120 89.820 ;
  LAYER ME2 ;
  RECT 0.000 86.580 1.120 89.820 ;
  LAYER ME1 ;
  RECT 0.000 86.580 1.120 89.820 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 47.380 1.120 50.620 ;
  LAYER ME3 ;
  RECT 0.000 47.380 1.120 50.620 ;
  LAYER ME2 ;
  RECT 0.000 47.380 1.120 50.620 ;
  LAYER ME1 ;
  RECT 0.000 47.380 1.120 50.620 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 39.540 1.120 42.780 ;
  LAYER ME3 ;
  RECT 0.000 39.540 1.120 42.780 ;
  LAYER ME2 ;
  RECT 0.000 39.540 1.120 42.780 ;
  LAYER ME1 ;
  RECT 0.000 39.540 1.120 42.780 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 31.700 1.120 34.940 ;
  LAYER ME3 ;
  RECT 0.000 31.700 1.120 34.940 ;
  LAYER ME2 ;
  RECT 0.000 31.700 1.120 34.940 ;
  LAYER ME1 ;
  RECT 0.000 31.700 1.120 34.940 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 23.860 1.120 27.100 ;
  LAYER ME3 ;
  RECT 0.000 23.860 1.120 27.100 ;
  LAYER ME2 ;
  RECT 0.000 23.860 1.120 27.100 ;
  LAYER ME1 ;
  RECT 0.000 23.860 1.120 27.100 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 16.020 1.120 19.260 ;
  LAYER ME3 ;
  RECT 0.000 16.020 1.120 19.260 ;
  LAYER ME2 ;
  RECT 0.000 16.020 1.120 19.260 ;
  LAYER ME1 ;
  RECT 0.000 16.020 1.120 19.260 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 8.180 1.120 11.420 ;
  LAYER ME3 ;
  RECT 0.000 8.180 1.120 11.420 ;
  LAYER ME2 ;
  RECT 0.000 8.180 1.120 11.420 ;
  LAYER ME1 ;
  RECT 0.000 8.180 1.120 11.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 980.000 175.280 983.540 176.400 ;
  LAYER ME3 ;
  RECT 980.000 175.280 983.540 176.400 ;
  LAYER ME2 ;
  RECT 980.000 175.280 983.540 176.400 ;
  LAYER ME1 ;
  RECT 980.000 175.280 983.540 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 971.320 175.280 974.860 176.400 ;
  LAYER ME3 ;
  RECT 971.320 175.280 974.860 176.400 ;
  LAYER ME2 ;
  RECT 971.320 175.280 974.860 176.400 ;
  LAYER ME1 ;
  RECT 971.320 175.280 974.860 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 962.640 175.280 966.180 176.400 ;
  LAYER ME3 ;
  RECT 962.640 175.280 966.180 176.400 ;
  LAYER ME2 ;
  RECT 962.640 175.280 966.180 176.400 ;
  LAYER ME1 ;
  RECT 962.640 175.280 966.180 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 919.240 175.280 922.780 176.400 ;
  LAYER ME3 ;
  RECT 919.240 175.280 922.780 176.400 ;
  LAYER ME2 ;
  RECT 919.240 175.280 922.780 176.400 ;
  LAYER ME1 ;
  RECT 919.240 175.280 922.780 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 910.560 175.280 914.100 176.400 ;
  LAYER ME3 ;
  RECT 910.560 175.280 914.100 176.400 ;
  LAYER ME2 ;
  RECT 910.560 175.280 914.100 176.400 ;
  LAYER ME1 ;
  RECT 910.560 175.280 914.100 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 901.880 175.280 905.420 176.400 ;
  LAYER ME3 ;
  RECT 901.880 175.280 905.420 176.400 ;
  LAYER ME2 ;
  RECT 901.880 175.280 905.420 176.400 ;
  LAYER ME1 ;
  RECT 901.880 175.280 905.420 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 893.200 175.280 896.740 176.400 ;
  LAYER ME3 ;
  RECT 893.200 175.280 896.740 176.400 ;
  LAYER ME2 ;
  RECT 893.200 175.280 896.740 176.400 ;
  LAYER ME1 ;
  RECT 893.200 175.280 896.740 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 884.520 175.280 888.060 176.400 ;
  LAYER ME3 ;
  RECT 884.520 175.280 888.060 176.400 ;
  LAYER ME2 ;
  RECT 884.520 175.280 888.060 176.400 ;
  LAYER ME1 ;
  RECT 884.520 175.280 888.060 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 875.840 175.280 879.380 176.400 ;
  LAYER ME3 ;
  RECT 875.840 175.280 879.380 176.400 ;
  LAYER ME2 ;
  RECT 875.840 175.280 879.380 176.400 ;
  LAYER ME1 ;
  RECT 875.840 175.280 879.380 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 832.440 175.280 835.980 176.400 ;
  LAYER ME3 ;
  RECT 832.440 175.280 835.980 176.400 ;
  LAYER ME2 ;
  RECT 832.440 175.280 835.980 176.400 ;
  LAYER ME1 ;
  RECT 832.440 175.280 835.980 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 823.760 175.280 827.300 176.400 ;
  LAYER ME3 ;
  RECT 823.760 175.280 827.300 176.400 ;
  LAYER ME2 ;
  RECT 823.760 175.280 827.300 176.400 ;
  LAYER ME1 ;
  RECT 823.760 175.280 827.300 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 815.080 175.280 818.620 176.400 ;
  LAYER ME3 ;
  RECT 815.080 175.280 818.620 176.400 ;
  LAYER ME2 ;
  RECT 815.080 175.280 818.620 176.400 ;
  LAYER ME1 ;
  RECT 815.080 175.280 818.620 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 806.400 175.280 809.940 176.400 ;
  LAYER ME3 ;
  RECT 806.400 175.280 809.940 176.400 ;
  LAYER ME2 ;
  RECT 806.400 175.280 809.940 176.400 ;
  LAYER ME1 ;
  RECT 806.400 175.280 809.940 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 797.720 175.280 801.260 176.400 ;
  LAYER ME3 ;
  RECT 797.720 175.280 801.260 176.400 ;
  LAYER ME2 ;
  RECT 797.720 175.280 801.260 176.400 ;
  LAYER ME1 ;
  RECT 797.720 175.280 801.260 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 789.040 175.280 792.580 176.400 ;
  LAYER ME3 ;
  RECT 789.040 175.280 792.580 176.400 ;
  LAYER ME2 ;
  RECT 789.040 175.280 792.580 176.400 ;
  LAYER ME1 ;
  RECT 789.040 175.280 792.580 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 745.640 175.280 749.180 176.400 ;
  LAYER ME3 ;
  RECT 745.640 175.280 749.180 176.400 ;
  LAYER ME2 ;
  RECT 745.640 175.280 749.180 176.400 ;
  LAYER ME1 ;
  RECT 745.640 175.280 749.180 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 736.960 175.280 740.500 176.400 ;
  LAYER ME3 ;
  RECT 736.960 175.280 740.500 176.400 ;
  LAYER ME2 ;
  RECT 736.960 175.280 740.500 176.400 ;
  LAYER ME1 ;
  RECT 736.960 175.280 740.500 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 728.280 175.280 731.820 176.400 ;
  LAYER ME3 ;
  RECT 728.280 175.280 731.820 176.400 ;
  LAYER ME2 ;
  RECT 728.280 175.280 731.820 176.400 ;
  LAYER ME1 ;
  RECT 728.280 175.280 731.820 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 719.600 175.280 723.140 176.400 ;
  LAYER ME3 ;
  RECT 719.600 175.280 723.140 176.400 ;
  LAYER ME2 ;
  RECT 719.600 175.280 723.140 176.400 ;
  LAYER ME1 ;
  RECT 719.600 175.280 723.140 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 710.920 175.280 714.460 176.400 ;
  LAYER ME3 ;
  RECT 710.920 175.280 714.460 176.400 ;
  LAYER ME2 ;
  RECT 710.920 175.280 714.460 176.400 ;
  LAYER ME1 ;
  RECT 710.920 175.280 714.460 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 702.240 175.280 705.780 176.400 ;
  LAYER ME3 ;
  RECT 702.240 175.280 705.780 176.400 ;
  LAYER ME2 ;
  RECT 702.240 175.280 705.780 176.400 ;
  LAYER ME1 ;
  RECT 702.240 175.280 705.780 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 658.840 175.280 662.380 176.400 ;
  LAYER ME3 ;
  RECT 658.840 175.280 662.380 176.400 ;
  LAYER ME2 ;
  RECT 658.840 175.280 662.380 176.400 ;
  LAYER ME1 ;
  RECT 658.840 175.280 662.380 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 650.160 175.280 653.700 176.400 ;
  LAYER ME3 ;
  RECT 650.160 175.280 653.700 176.400 ;
  LAYER ME2 ;
  RECT 650.160 175.280 653.700 176.400 ;
  LAYER ME1 ;
  RECT 650.160 175.280 653.700 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 641.480 175.280 645.020 176.400 ;
  LAYER ME3 ;
  RECT 641.480 175.280 645.020 176.400 ;
  LAYER ME2 ;
  RECT 641.480 175.280 645.020 176.400 ;
  LAYER ME1 ;
  RECT 641.480 175.280 645.020 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 632.800 175.280 636.340 176.400 ;
  LAYER ME3 ;
  RECT 632.800 175.280 636.340 176.400 ;
  LAYER ME2 ;
  RECT 632.800 175.280 636.340 176.400 ;
  LAYER ME1 ;
  RECT 632.800 175.280 636.340 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 624.120 175.280 627.660 176.400 ;
  LAYER ME3 ;
  RECT 624.120 175.280 627.660 176.400 ;
  LAYER ME2 ;
  RECT 624.120 175.280 627.660 176.400 ;
  LAYER ME1 ;
  RECT 624.120 175.280 627.660 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 615.440 175.280 618.980 176.400 ;
  LAYER ME3 ;
  RECT 615.440 175.280 618.980 176.400 ;
  LAYER ME2 ;
  RECT 615.440 175.280 618.980 176.400 ;
  LAYER ME1 ;
  RECT 615.440 175.280 618.980 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 572.040 175.280 575.580 176.400 ;
  LAYER ME3 ;
  RECT 572.040 175.280 575.580 176.400 ;
  LAYER ME2 ;
  RECT 572.040 175.280 575.580 176.400 ;
  LAYER ME1 ;
  RECT 572.040 175.280 575.580 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 563.360 175.280 566.900 176.400 ;
  LAYER ME3 ;
  RECT 563.360 175.280 566.900 176.400 ;
  LAYER ME2 ;
  RECT 563.360 175.280 566.900 176.400 ;
  LAYER ME1 ;
  RECT 563.360 175.280 566.900 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 554.680 175.280 558.220 176.400 ;
  LAYER ME3 ;
  RECT 554.680 175.280 558.220 176.400 ;
  LAYER ME2 ;
  RECT 554.680 175.280 558.220 176.400 ;
  LAYER ME1 ;
  RECT 554.680 175.280 558.220 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 546.000 175.280 549.540 176.400 ;
  LAYER ME3 ;
  RECT 546.000 175.280 549.540 176.400 ;
  LAYER ME2 ;
  RECT 546.000 175.280 549.540 176.400 ;
  LAYER ME1 ;
  RECT 546.000 175.280 549.540 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 537.320 175.280 540.860 176.400 ;
  LAYER ME3 ;
  RECT 537.320 175.280 540.860 176.400 ;
  LAYER ME2 ;
  RECT 537.320 175.280 540.860 176.400 ;
  LAYER ME1 ;
  RECT 537.320 175.280 540.860 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 528.640 175.280 532.180 176.400 ;
  LAYER ME3 ;
  RECT 528.640 175.280 532.180 176.400 ;
  LAYER ME2 ;
  RECT 528.640 175.280 532.180 176.400 ;
  LAYER ME1 ;
  RECT 528.640 175.280 532.180 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 485.240 175.280 488.780 176.400 ;
  LAYER ME3 ;
  RECT 485.240 175.280 488.780 176.400 ;
  LAYER ME2 ;
  RECT 485.240 175.280 488.780 176.400 ;
  LAYER ME1 ;
  RECT 485.240 175.280 488.780 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 476.560 175.280 480.100 176.400 ;
  LAYER ME3 ;
  RECT 476.560 175.280 480.100 176.400 ;
  LAYER ME2 ;
  RECT 476.560 175.280 480.100 176.400 ;
  LAYER ME1 ;
  RECT 476.560 175.280 480.100 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 467.880 175.280 471.420 176.400 ;
  LAYER ME3 ;
  RECT 467.880 175.280 471.420 176.400 ;
  LAYER ME2 ;
  RECT 467.880 175.280 471.420 176.400 ;
  LAYER ME1 ;
  RECT 467.880 175.280 471.420 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 459.200 175.280 462.740 176.400 ;
  LAYER ME3 ;
  RECT 459.200 175.280 462.740 176.400 ;
  LAYER ME2 ;
  RECT 459.200 175.280 462.740 176.400 ;
  LAYER ME1 ;
  RECT 459.200 175.280 462.740 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 450.520 175.280 454.060 176.400 ;
  LAYER ME3 ;
  RECT 450.520 175.280 454.060 176.400 ;
  LAYER ME2 ;
  RECT 450.520 175.280 454.060 176.400 ;
  LAYER ME1 ;
  RECT 450.520 175.280 454.060 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 441.840 175.280 445.380 176.400 ;
  LAYER ME3 ;
  RECT 441.840 175.280 445.380 176.400 ;
  LAYER ME2 ;
  RECT 441.840 175.280 445.380 176.400 ;
  LAYER ME1 ;
  RECT 441.840 175.280 445.380 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 398.440 175.280 401.980 176.400 ;
  LAYER ME3 ;
  RECT 398.440 175.280 401.980 176.400 ;
  LAYER ME2 ;
  RECT 398.440 175.280 401.980 176.400 ;
  LAYER ME1 ;
  RECT 398.440 175.280 401.980 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 389.760 175.280 393.300 176.400 ;
  LAYER ME3 ;
  RECT 389.760 175.280 393.300 176.400 ;
  LAYER ME2 ;
  RECT 389.760 175.280 393.300 176.400 ;
  LAYER ME1 ;
  RECT 389.760 175.280 393.300 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 381.080 175.280 384.620 176.400 ;
  LAYER ME3 ;
  RECT 381.080 175.280 384.620 176.400 ;
  LAYER ME2 ;
  RECT 381.080 175.280 384.620 176.400 ;
  LAYER ME1 ;
  RECT 381.080 175.280 384.620 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 372.400 175.280 375.940 176.400 ;
  LAYER ME3 ;
  RECT 372.400 175.280 375.940 176.400 ;
  LAYER ME2 ;
  RECT 372.400 175.280 375.940 176.400 ;
  LAYER ME1 ;
  RECT 372.400 175.280 375.940 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 363.720 175.280 367.260 176.400 ;
  LAYER ME3 ;
  RECT 363.720 175.280 367.260 176.400 ;
  LAYER ME2 ;
  RECT 363.720 175.280 367.260 176.400 ;
  LAYER ME1 ;
  RECT 363.720 175.280 367.260 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 355.040 175.280 358.580 176.400 ;
  LAYER ME3 ;
  RECT 355.040 175.280 358.580 176.400 ;
  LAYER ME2 ;
  RECT 355.040 175.280 358.580 176.400 ;
  LAYER ME1 ;
  RECT 355.040 175.280 358.580 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 311.640 175.280 315.180 176.400 ;
  LAYER ME3 ;
  RECT 311.640 175.280 315.180 176.400 ;
  LAYER ME2 ;
  RECT 311.640 175.280 315.180 176.400 ;
  LAYER ME1 ;
  RECT 311.640 175.280 315.180 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 302.960 175.280 306.500 176.400 ;
  LAYER ME3 ;
  RECT 302.960 175.280 306.500 176.400 ;
  LAYER ME2 ;
  RECT 302.960 175.280 306.500 176.400 ;
  LAYER ME1 ;
  RECT 302.960 175.280 306.500 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 294.280 175.280 297.820 176.400 ;
  LAYER ME3 ;
  RECT 294.280 175.280 297.820 176.400 ;
  LAYER ME2 ;
  RECT 294.280 175.280 297.820 176.400 ;
  LAYER ME1 ;
  RECT 294.280 175.280 297.820 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 285.600 175.280 289.140 176.400 ;
  LAYER ME3 ;
  RECT 285.600 175.280 289.140 176.400 ;
  LAYER ME2 ;
  RECT 285.600 175.280 289.140 176.400 ;
  LAYER ME1 ;
  RECT 285.600 175.280 289.140 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 276.920 175.280 280.460 176.400 ;
  LAYER ME3 ;
  RECT 276.920 175.280 280.460 176.400 ;
  LAYER ME2 ;
  RECT 276.920 175.280 280.460 176.400 ;
  LAYER ME1 ;
  RECT 276.920 175.280 280.460 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 268.240 175.280 271.780 176.400 ;
  LAYER ME3 ;
  RECT 268.240 175.280 271.780 176.400 ;
  LAYER ME2 ;
  RECT 268.240 175.280 271.780 176.400 ;
  LAYER ME1 ;
  RECT 268.240 175.280 271.780 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 224.840 175.280 228.380 176.400 ;
  LAYER ME3 ;
  RECT 224.840 175.280 228.380 176.400 ;
  LAYER ME2 ;
  RECT 224.840 175.280 228.380 176.400 ;
  LAYER ME1 ;
  RECT 224.840 175.280 228.380 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 216.160 175.280 219.700 176.400 ;
  LAYER ME3 ;
  RECT 216.160 175.280 219.700 176.400 ;
  LAYER ME2 ;
  RECT 216.160 175.280 219.700 176.400 ;
  LAYER ME1 ;
  RECT 216.160 175.280 219.700 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 207.480 175.280 211.020 176.400 ;
  LAYER ME3 ;
  RECT 207.480 175.280 211.020 176.400 ;
  LAYER ME2 ;
  RECT 207.480 175.280 211.020 176.400 ;
  LAYER ME1 ;
  RECT 207.480 175.280 211.020 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 198.800 175.280 202.340 176.400 ;
  LAYER ME3 ;
  RECT 198.800 175.280 202.340 176.400 ;
  LAYER ME2 ;
  RECT 198.800 175.280 202.340 176.400 ;
  LAYER ME1 ;
  RECT 198.800 175.280 202.340 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 190.120 175.280 193.660 176.400 ;
  LAYER ME3 ;
  RECT 190.120 175.280 193.660 176.400 ;
  LAYER ME2 ;
  RECT 190.120 175.280 193.660 176.400 ;
  LAYER ME1 ;
  RECT 190.120 175.280 193.660 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 181.440 175.280 184.980 176.400 ;
  LAYER ME3 ;
  RECT 181.440 175.280 184.980 176.400 ;
  LAYER ME2 ;
  RECT 181.440 175.280 184.980 176.400 ;
  LAYER ME1 ;
  RECT 181.440 175.280 184.980 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 138.040 175.280 141.580 176.400 ;
  LAYER ME3 ;
  RECT 138.040 175.280 141.580 176.400 ;
  LAYER ME2 ;
  RECT 138.040 175.280 141.580 176.400 ;
  LAYER ME1 ;
  RECT 138.040 175.280 141.580 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 129.360 175.280 132.900 176.400 ;
  LAYER ME3 ;
  RECT 129.360 175.280 132.900 176.400 ;
  LAYER ME2 ;
  RECT 129.360 175.280 132.900 176.400 ;
  LAYER ME1 ;
  RECT 129.360 175.280 132.900 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 120.680 175.280 124.220 176.400 ;
  LAYER ME3 ;
  RECT 120.680 175.280 124.220 176.400 ;
  LAYER ME2 ;
  RECT 120.680 175.280 124.220 176.400 ;
  LAYER ME1 ;
  RECT 120.680 175.280 124.220 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 112.000 175.280 115.540 176.400 ;
  LAYER ME3 ;
  RECT 112.000 175.280 115.540 176.400 ;
  LAYER ME2 ;
  RECT 112.000 175.280 115.540 176.400 ;
  LAYER ME1 ;
  RECT 112.000 175.280 115.540 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 103.320 175.280 106.860 176.400 ;
  LAYER ME3 ;
  RECT 103.320 175.280 106.860 176.400 ;
  LAYER ME2 ;
  RECT 103.320 175.280 106.860 176.400 ;
  LAYER ME1 ;
  RECT 103.320 175.280 106.860 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 94.640 175.280 98.180 176.400 ;
  LAYER ME3 ;
  RECT 94.640 175.280 98.180 176.400 ;
  LAYER ME2 ;
  RECT 94.640 175.280 98.180 176.400 ;
  LAYER ME1 ;
  RECT 94.640 175.280 98.180 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 51.240 175.280 54.780 176.400 ;
  LAYER ME3 ;
  RECT 51.240 175.280 54.780 176.400 ;
  LAYER ME2 ;
  RECT 51.240 175.280 54.780 176.400 ;
  LAYER ME1 ;
  RECT 51.240 175.280 54.780 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 42.560 175.280 46.100 176.400 ;
  LAYER ME3 ;
  RECT 42.560 175.280 46.100 176.400 ;
  LAYER ME2 ;
  RECT 42.560 175.280 46.100 176.400 ;
  LAYER ME1 ;
  RECT 42.560 175.280 46.100 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 33.880 175.280 37.420 176.400 ;
  LAYER ME3 ;
  RECT 33.880 175.280 37.420 176.400 ;
  LAYER ME2 ;
  RECT 33.880 175.280 37.420 176.400 ;
  LAYER ME1 ;
  RECT 33.880 175.280 37.420 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 25.200 175.280 28.740 176.400 ;
  LAYER ME3 ;
  RECT 25.200 175.280 28.740 176.400 ;
  LAYER ME2 ;
  RECT 25.200 175.280 28.740 176.400 ;
  LAYER ME1 ;
  RECT 25.200 175.280 28.740 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 16.520 175.280 20.060 176.400 ;
  LAYER ME3 ;
  RECT 16.520 175.280 20.060 176.400 ;
  LAYER ME2 ;
  RECT 16.520 175.280 20.060 176.400 ;
  LAYER ME1 ;
  RECT 16.520 175.280 20.060 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 7.840 175.280 11.380 176.400 ;
  LAYER ME3 ;
  RECT 7.840 175.280 11.380 176.400 ;
  LAYER ME2 ;
  RECT 7.840 175.280 11.380 176.400 ;
  LAYER ME1 ;
  RECT 7.840 175.280 11.380 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 983.100 0.000 986.640 1.120 ;
  LAYER ME3 ;
  RECT 983.100 0.000 986.640 1.120 ;
  LAYER ME2 ;
  RECT 983.100 0.000 986.640 1.120 ;
  LAYER ME1 ;
  RECT 983.100 0.000 986.640 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 961.400 0.000 964.940 1.120 ;
  LAYER ME3 ;
  RECT 961.400 0.000 964.940 1.120 ;
  LAYER ME2 ;
  RECT 961.400 0.000 964.940 1.120 ;
  LAYER ME1 ;
  RECT 961.400 0.000 964.940 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 944.660 0.000 948.200 1.120 ;
  LAYER ME3 ;
  RECT 944.660 0.000 948.200 1.120 ;
  LAYER ME2 ;
  RECT 944.660 0.000 948.200 1.120 ;
  LAYER ME1 ;
  RECT 944.660 0.000 948.200 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 918.000 0.000 921.540 1.120 ;
  LAYER ME3 ;
  RECT 918.000 0.000 921.540 1.120 ;
  LAYER ME2 ;
  RECT 918.000 0.000 921.540 1.120 ;
  LAYER ME1 ;
  RECT 918.000 0.000 921.540 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 896.920 0.000 900.460 1.120 ;
  LAYER ME3 ;
  RECT 896.920 0.000 900.460 1.120 ;
  LAYER ME2 ;
  RECT 896.920 0.000 900.460 1.120 ;
  LAYER ME1 ;
  RECT 896.920 0.000 900.460 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 783.460 0.000 787.000 1.120 ;
  LAYER ME3 ;
  RECT 783.460 0.000 787.000 1.120 ;
  LAYER ME2 ;
  RECT 783.460 0.000 787.000 1.120 ;
  LAYER ME1 ;
  RECT 783.460 0.000 787.000 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 761.760 0.000 765.300 1.120 ;
  LAYER ME3 ;
  RECT 761.760 0.000 765.300 1.120 ;
  LAYER ME2 ;
  RECT 761.760 0.000 765.300 1.120 ;
  LAYER ME1 ;
  RECT 761.760 0.000 765.300 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 735.100 0.000 738.640 1.120 ;
  LAYER ME3 ;
  RECT 735.100 0.000 738.640 1.120 ;
  LAYER ME2 ;
  RECT 735.100 0.000 738.640 1.120 ;
  LAYER ME1 ;
  RECT 735.100 0.000 738.640 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 718.980 0.000 722.520 1.120 ;
  LAYER ME3 ;
  RECT 718.980 0.000 722.520 1.120 ;
  LAYER ME2 ;
  RECT 718.980 0.000 722.520 1.120 ;
  LAYER ME1 ;
  RECT 718.980 0.000 722.520 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 692.320 0.000 695.860 1.120 ;
  LAYER ME3 ;
  RECT 692.320 0.000 695.860 1.120 ;
  LAYER ME2 ;
  RECT 692.320 0.000 695.860 1.120 ;
  LAYER ME1 ;
  RECT 692.320 0.000 695.860 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 670.620 0.000 674.160 1.120 ;
  LAYER ME3 ;
  RECT 670.620 0.000 674.160 1.120 ;
  LAYER ME2 ;
  RECT 670.620 0.000 674.160 1.120 ;
  LAYER ME1 ;
  RECT 670.620 0.000 674.160 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 557.780 0.000 561.320 1.120 ;
  LAYER ME3 ;
  RECT 557.780 0.000 561.320 1.120 ;
  LAYER ME2 ;
  RECT 557.780 0.000 561.320 1.120 ;
  LAYER ME1 ;
  RECT 557.780 0.000 561.320 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 536.080 0.000 539.620 1.120 ;
  LAYER ME3 ;
  RECT 536.080 0.000 539.620 1.120 ;
  LAYER ME2 ;
  RECT 536.080 0.000 539.620 1.120 ;
  LAYER ME1 ;
  RECT 536.080 0.000 539.620 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 508.800 0.000 512.340 1.120 ;
  LAYER ME3 ;
  RECT 508.800 0.000 512.340 1.120 ;
  LAYER ME2 ;
  RECT 508.800 0.000 512.340 1.120 ;
  LAYER ME1 ;
  RECT 508.800 0.000 512.340 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 500.120 0.000 503.660 1.120 ;
  LAYER ME3 ;
  RECT 500.120 0.000 503.660 1.120 ;
  LAYER ME2 ;
  RECT 500.120 0.000 503.660 1.120 ;
  LAYER ME1 ;
  RECT 500.120 0.000 503.660 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 472.220 0.000 475.760 1.120 ;
  LAYER ME3 ;
  RECT 472.220 0.000 475.760 1.120 ;
  LAYER ME2 ;
  RECT 472.220 0.000 475.760 1.120 ;
  LAYER ME1 ;
  RECT 472.220 0.000 475.760 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 461.060 0.000 464.600 1.120 ;
  LAYER ME3 ;
  RECT 461.060 0.000 464.600 1.120 ;
  LAYER ME2 ;
  RECT 461.060 0.000 464.600 1.120 ;
  LAYER ME1 ;
  RECT 461.060 0.000 464.600 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 353.180 0.000 356.720 1.120 ;
  LAYER ME3 ;
  RECT 353.180 0.000 356.720 1.120 ;
  LAYER ME2 ;
  RECT 353.180 0.000 356.720 1.120 ;
  LAYER ME1 ;
  RECT 353.180 0.000 356.720 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 326.520 0.000 330.060 1.120 ;
  LAYER ME3 ;
  RECT 326.520 0.000 330.060 1.120 ;
  LAYER ME2 ;
  RECT 326.520 0.000 330.060 1.120 ;
  LAYER ME1 ;
  RECT 326.520 0.000 330.060 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 309.780 0.000 313.320 1.120 ;
  LAYER ME3 ;
  RECT 309.780 0.000 313.320 1.120 ;
  LAYER ME2 ;
  RECT 309.780 0.000 313.320 1.120 ;
  LAYER ME1 ;
  RECT 309.780 0.000 313.320 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 283.120 0.000 286.660 1.120 ;
  LAYER ME3 ;
  RECT 283.120 0.000 286.660 1.120 ;
  LAYER ME2 ;
  RECT 283.120 0.000 286.660 1.120 ;
  LAYER ME1 ;
  RECT 283.120 0.000 286.660 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 261.420 0.000 264.960 1.120 ;
  LAYER ME3 ;
  RECT 261.420 0.000 264.960 1.120 ;
  LAYER ME2 ;
  RECT 261.420 0.000 264.960 1.120 ;
  LAYER ME1 ;
  RECT 261.420 0.000 264.960 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 239.720 0.000 243.260 1.120 ;
  LAYER ME3 ;
  RECT 239.720 0.000 243.260 1.120 ;
  LAYER ME2 ;
  RECT 239.720 0.000 243.260 1.120 ;
  LAYER ME1 ;
  RECT 239.720 0.000 243.260 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 126.880 0.000 130.420 1.120 ;
  LAYER ME3 ;
  RECT 126.880 0.000 130.420 1.120 ;
  LAYER ME2 ;
  RECT 126.880 0.000 130.420 1.120 ;
  LAYER ME1 ;
  RECT 126.880 0.000 130.420 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 100.220 0.000 103.760 1.120 ;
  LAYER ME3 ;
  RECT 100.220 0.000 103.760 1.120 ;
  LAYER ME2 ;
  RECT 100.220 0.000 103.760 1.120 ;
  LAYER ME1 ;
  RECT 100.220 0.000 103.760 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 83.480 0.000 87.020 1.120 ;
  LAYER ME3 ;
  RECT 83.480 0.000 87.020 1.120 ;
  LAYER ME2 ;
  RECT 83.480 0.000 87.020 1.120 ;
  LAYER ME1 ;
  RECT 83.480 0.000 87.020 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 56.820 0.000 60.360 1.120 ;
  LAYER ME3 ;
  RECT 56.820 0.000 60.360 1.120 ;
  LAYER ME2 ;
  RECT 56.820 0.000 60.360 1.120 ;
  LAYER ME1 ;
  RECT 56.820 0.000 60.360 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 35.740 0.000 39.280 1.120 ;
  LAYER ME3 ;
  RECT 35.740 0.000 39.280 1.120 ;
  LAYER ME2 ;
  RECT 35.740 0.000 39.280 1.120 ;
  LAYER ME1 ;
  RECT 35.740 0.000 39.280 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 14.040 0.000 17.580 1.120 ;
  LAYER ME3 ;
  RECT 14.040 0.000 17.580 1.120 ;
  LAYER ME2 ;
  RECT 14.040 0.000 17.580 1.120 ;
  LAYER ME1 ;
  RECT 14.040 0.000 17.580 1.120 ;
 END
END VCC
PIN GND
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
 PORT
  LAYER ME4 ;
  RECT 993.360 129.700 994.480 132.940 ;
  LAYER ME3 ;
  RECT 993.360 129.700 994.480 132.940 ;
  LAYER ME2 ;
  RECT 993.360 129.700 994.480 132.940 ;
  LAYER ME1 ;
  RECT 993.360 129.700 994.480 132.940 ;
 END
 PORT
  LAYER ME4 ;
  RECT 993.360 121.860 994.480 125.100 ;
  LAYER ME3 ;
  RECT 993.360 121.860 994.480 125.100 ;
  LAYER ME2 ;
  RECT 993.360 121.860 994.480 125.100 ;
  LAYER ME1 ;
  RECT 993.360 121.860 994.480 125.100 ;
 END
 PORT
  LAYER ME4 ;
  RECT 993.360 114.020 994.480 117.260 ;
  LAYER ME3 ;
  RECT 993.360 114.020 994.480 117.260 ;
  LAYER ME2 ;
  RECT 993.360 114.020 994.480 117.260 ;
  LAYER ME1 ;
  RECT 993.360 114.020 994.480 117.260 ;
 END
 PORT
  LAYER ME4 ;
  RECT 993.360 106.180 994.480 109.420 ;
  LAYER ME3 ;
  RECT 993.360 106.180 994.480 109.420 ;
  LAYER ME2 ;
  RECT 993.360 106.180 994.480 109.420 ;
  LAYER ME1 ;
  RECT 993.360 106.180 994.480 109.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 993.360 98.340 994.480 101.580 ;
  LAYER ME3 ;
  RECT 993.360 98.340 994.480 101.580 ;
  LAYER ME2 ;
  RECT 993.360 98.340 994.480 101.580 ;
  LAYER ME1 ;
  RECT 993.360 98.340 994.480 101.580 ;
 END
 PORT
  LAYER ME4 ;
  RECT 993.360 90.500 994.480 93.740 ;
  LAYER ME3 ;
  RECT 993.360 90.500 994.480 93.740 ;
  LAYER ME2 ;
  RECT 993.360 90.500 994.480 93.740 ;
  LAYER ME1 ;
  RECT 993.360 90.500 994.480 93.740 ;
 END
 PORT
  LAYER ME4 ;
  RECT 993.360 51.300 994.480 54.540 ;
  LAYER ME3 ;
  RECT 993.360 51.300 994.480 54.540 ;
  LAYER ME2 ;
  RECT 993.360 51.300 994.480 54.540 ;
  LAYER ME1 ;
  RECT 993.360 51.300 994.480 54.540 ;
 END
 PORT
  LAYER ME4 ;
  RECT 993.360 43.460 994.480 46.700 ;
  LAYER ME3 ;
  RECT 993.360 43.460 994.480 46.700 ;
  LAYER ME2 ;
  RECT 993.360 43.460 994.480 46.700 ;
  LAYER ME1 ;
  RECT 993.360 43.460 994.480 46.700 ;
 END
 PORT
  LAYER ME4 ;
  RECT 993.360 35.620 994.480 38.860 ;
  LAYER ME3 ;
  RECT 993.360 35.620 994.480 38.860 ;
  LAYER ME2 ;
  RECT 993.360 35.620 994.480 38.860 ;
  LAYER ME1 ;
  RECT 993.360 35.620 994.480 38.860 ;
 END
 PORT
  LAYER ME4 ;
  RECT 993.360 27.780 994.480 31.020 ;
  LAYER ME3 ;
  RECT 993.360 27.780 994.480 31.020 ;
  LAYER ME2 ;
  RECT 993.360 27.780 994.480 31.020 ;
  LAYER ME1 ;
  RECT 993.360 27.780 994.480 31.020 ;
 END
 PORT
  LAYER ME4 ;
  RECT 993.360 19.940 994.480 23.180 ;
  LAYER ME3 ;
  RECT 993.360 19.940 994.480 23.180 ;
  LAYER ME2 ;
  RECT 993.360 19.940 994.480 23.180 ;
  LAYER ME1 ;
  RECT 993.360 19.940 994.480 23.180 ;
 END
 PORT
  LAYER ME4 ;
  RECT 993.360 12.100 994.480 15.340 ;
  LAYER ME3 ;
  RECT 993.360 12.100 994.480 15.340 ;
  LAYER ME2 ;
  RECT 993.360 12.100 994.480 15.340 ;
  LAYER ME1 ;
  RECT 993.360 12.100 994.480 15.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 129.700 1.120 132.940 ;
  LAYER ME3 ;
  RECT 0.000 129.700 1.120 132.940 ;
  LAYER ME2 ;
  RECT 0.000 129.700 1.120 132.940 ;
  LAYER ME1 ;
  RECT 0.000 129.700 1.120 132.940 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 121.860 1.120 125.100 ;
  LAYER ME3 ;
  RECT 0.000 121.860 1.120 125.100 ;
  LAYER ME2 ;
  RECT 0.000 121.860 1.120 125.100 ;
  LAYER ME1 ;
  RECT 0.000 121.860 1.120 125.100 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 114.020 1.120 117.260 ;
  LAYER ME3 ;
  RECT 0.000 114.020 1.120 117.260 ;
  LAYER ME2 ;
  RECT 0.000 114.020 1.120 117.260 ;
  LAYER ME1 ;
  RECT 0.000 114.020 1.120 117.260 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 106.180 1.120 109.420 ;
  LAYER ME3 ;
  RECT 0.000 106.180 1.120 109.420 ;
  LAYER ME2 ;
  RECT 0.000 106.180 1.120 109.420 ;
  LAYER ME1 ;
  RECT 0.000 106.180 1.120 109.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 98.340 1.120 101.580 ;
  LAYER ME3 ;
  RECT 0.000 98.340 1.120 101.580 ;
  LAYER ME2 ;
  RECT 0.000 98.340 1.120 101.580 ;
  LAYER ME1 ;
  RECT 0.000 98.340 1.120 101.580 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 90.500 1.120 93.740 ;
  LAYER ME3 ;
  RECT 0.000 90.500 1.120 93.740 ;
  LAYER ME2 ;
  RECT 0.000 90.500 1.120 93.740 ;
  LAYER ME1 ;
  RECT 0.000 90.500 1.120 93.740 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 51.300 1.120 54.540 ;
  LAYER ME3 ;
  RECT 0.000 51.300 1.120 54.540 ;
  LAYER ME2 ;
  RECT 0.000 51.300 1.120 54.540 ;
  LAYER ME1 ;
  RECT 0.000 51.300 1.120 54.540 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 43.460 1.120 46.700 ;
  LAYER ME3 ;
  RECT 0.000 43.460 1.120 46.700 ;
  LAYER ME2 ;
  RECT 0.000 43.460 1.120 46.700 ;
  LAYER ME1 ;
  RECT 0.000 43.460 1.120 46.700 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 35.620 1.120 38.860 ;
  LAYER ME3 ;
  RECT 0.000 35.620 1.120 38.860 ;
  LAYER ME2 ;
  RECT 0.000 35.620 1.120 38.860 ;
  LAYER ME1 ;
  RECT 0.000 35.620 1.120 38.860 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 27.780 1.120 31.020 ;
  LAYER ME3 ;
  RECT 0.000 27.780 1.120 31.020 ;
  LAYER ME2 ;
  RECT 0.000 27.780 1.120 31.020 ;
  LAYER ME1 ;
  RECT 0.000 27.780 1.120 31.020 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 19.940 1.120 23.180 ;
  LAYER ME3 ;
  RECT 0.000 19.940 1.120 23.180 ;
  LAYER ME2 ;
  RECT 0.000 19.940 1.120 23.180 ;
  LAYER ME1 ;
  RECT 0.000 19.940 1.120 23.180 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 12.100 1.120 15.340 ;
  LAYER ME3 ;
  RECT 0.000 12.100 1.120 15.340 ;
  LAYER ME2 ;
  RECT 0.000 12.100 1.120 15.340 ;
  LAYER ME1 ;
  RECT 0.000 12.100 1.120 15.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 975.660 175.280 979.200 176.400 ;
  LAYER ME3 ;
  RECT 975.660 175.280 979.200 176.400 ;
  LAYER ME2 ;
  RECT 975.660 175.280 979.200 176.400 ;
  LAYER ME1 ;
  RECT 975.660 175.280 979.200 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 966.980 175.280 970.520 176.400 ;
  LAYER ME3 ;
  RECT 966.980 175.280 970.520 176.400 ;
  LAYER ME2 ;
  RECT 966.980 175.280 970.520 176.400 ;
  LAYER ME1 ;
  RECT 966.980 175.280 970.520 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 923.580 175.280 927.120 176.400 ;
  LAYER ME3 ;
  RECT 923.580 175.280 927.120 176.400 ;
  LAYER ME2 ;
  RECT 923.580 175.280 927.120 176.400 ;
  LAYER ME1 ;
  RECT 923.580 175.280 927.120 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 914.900 175.280 918.440 176.400 ;
  LAYER ME3 ;
  RECT 914.900 175.280 918.440 176.400 ;
  LAYER ME2 ;
  RECT 914.900 175.280 918.440 176.400 ;
  LAYER ME1 ;
  RECT 914.900 175.280 918.440 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 906.220 175.280 909.760 176.400 ;
  LAYER ME3 ;
  RECT 906.220 175.280 909.760 176.400 ;
  LAYER ME2 ;
  RECT 906.220 175.280 909.760 176.400 ;
  LAYER ME1 ;
  RECT 906.220 175.280 909.760 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 897.540 175.280 901.080 176.400 ;
  LAYER ME3 ;
  RECT 897.540 175.280 901.080 176.400 ;
  LAYER ME2 ;
  RECT 897.540 175.280 901.080 176.400 ;
  LAYER ME1 ;
  RECT 897.540 175.280 901.080 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 888.860 175.280 892.400 176.400 ;
  LAYER ME3 ;
  RECT 888.860 175.280 892.400 176.400 ;
  LAYER ME2 ;
  RECT 888.860 175.280 892.400 176.400 ;
  LAYER ME1 ;
  RECT 888.860 175.280 892.400 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 880.180 175.280 883.720 176.400 ;
  LAYER ME3 ;
  RECT 880.180 175.280 883.720 176.400 ;
  LAYER ME2 ;
  RECT 880.180 175.280 883.720 176.400 ;
  LAYER ME1 ;
  RECT 880.180 175.280 883.720 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 836.780 175.280 840.320 176.400 ;
  LAYER ME3 ;
  RECT 836.780 175.280 840.320 176.400 ;
  LAYER ME2 ;
  RECT 836.780 175.280 840.320 176.400 ;
  LAYER ME1 ;
  RECT 836.780 175.280 840.320 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 828.100 175.280 831.640 176.400 ;
  LAYER ME3 ;
  RECT 828.100 175.280 831.640 176.400 ;
  LAYER ME2 ;
  RECT 828.100 175.280 831.640 176.400 ;
  LAYER ME1 ;
  RECT 828.100 175.280 831.640 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 819.420 175.280 822.960 176.400 ;
  LAYER ME3 ;
  RECT 819.420 175.280 822.960 176.400 ;
  LAYER ME2 ;
  RECT 819.420 175.280 822.960 176.400 ;
  LAYER ME1 ;
  RECT 819.420 175.280 822.960 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 810.740 175.280 814.280 176.400 ;
  LAYER ME3 ;
  RECT 810.740 175.280 814.280 176.400 ;
  LAYER ME2 ;
  RECT 810.740 175.280 814.280 176.400 ;
  LAYER ME1 ;
  RECT 810.740 175.280 814.280 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 802.060 175.280 805.600 176.400 ;
  LAYER ME3 ;
  RECT 802.060 175.280 805.600 176.400 ;
  LAYER ME2 ;
  RECT 802.060 175.280 805.600 176.400 ;
  LAYER ME1 ;
  RECT 802.060 175.280 805.600 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 793.380 175.280 796.920 176.400 ;
  LAYER ME3 ;
  RECT 793.380 175.280 796.920 176.400 ;
  LAYER ME2 ;
  RECT 793.380 175.280 796.920 176.400 ;
  LAYER ME1 ;
  RECT 793.380 175.280 796.920 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 749.980 175.280 753.520 176.400 ;
  LAYER ME3 ;
  RECT 749.980 175.280 753.520 176.400 ;
  LAYER ME2 ;
  RECT 749.980 175.280 753.520 176.400 ;
  LAYER ME1 ;
  RECT 749.980 175.280 753.520 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 741.300 175.280 744.840 176.400 ;
  LAYER ME3 ;
  RECT 741.300 175.280 744.840 176.400 ;
  LAYER ME2 ;
  RECT 741.300 175.280 744.840 176.400 ;
  LAYER ME1 ;
  RECT 741.300 175.280 744.840 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 732.620 175.280 736.160 176.400 ;
  LAYER ME3 ;
  RECT 732.620 175.280 736.160 176.400 ;
  LAYER ME2 ;
  RECT 732.620 175.280 736.160 176.400 ;
  LAYER ME1 ;
  RECT 732.620 175.280 736.160 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 723.940 175.280 727.480 176.400 ;
  LAYER ME3 ;
  RECT 723.940 175.280 727.480 176.400 ;
  LAYER ME2 ;
  RECT 723.940 175.280 727.480 176.400 ;
  LAYER ME1 ;
  RECT 723.940 175.280 727.480 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 715.260 175.280 718.800 176.400 ;
  LAYER ME3 ;
  RECT 715.260 175.280 718.800 176.400 ;
  LAYER ME2 ;
  RECT 715.260 175.280 718.800 176.400 ;
  LAYER ME1 ;
  RECT 715.260 175.280 718.800 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 706.580 175.280 710.120 176.400 ;
  LAYER ME3 ;
  RECT 706.580 175.280 710.120 176.400 ;
  LAYER ME2 ;
  RECT 706.580 175.280 710.120 176.400 ;
  LAYER ME1 ;
  RECT 706.580 175.280 710.120 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 663.180 175.280 666.720 176.400 ;
  LAYER ME3 ;
  RECT 663.180 175.280 666.720 176.400 ;
  LAYER ME2 ;
  RECT 663.180 175.280 666.720 176.400 ;
  LAYER ME1 ;
  RECT 663.180 175.280 666.720 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 654.500 175.280 658.040 176.400 ;
  LAYER ME3 ;
  RECT 654.500 175.280 658.040 176.400 ;
  LAYER ME2 ;
  RECT 654.500 175.280 658.040 176.400 ;
  LAYER ME1 ;
  RECT 654.500 175.280 658.040 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 645.820 175.280 649.360 176.400 ;
  LAYER ME3 ;
  RECT 645.820 175.280 649.360 176.400 ;
  LAYER ME2 ;
  RECT 645.820 175.280 649.360 176.400 ;
  LAYER ME1 ;
  RECT 645.820 175.280 649.360 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 637.140 175.280 640.680 176.400 ;
  LAYER ME3 ;
  RECT 637.140 175.280 640.680 176.400 ;
  LAYER ME2 ;
  RECT 637.140 175.280 640.680 176.400 ;
  LAYER ME1 ;
  RECT 637.140 175.280 640.680 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 628.460 175.280 632.000 176.400 ;
  LAYER ME3 ;
  RECT 628.460 175.280 632.000 176.400 ;
  LAYER ME2 ;
  RECT 628.460 175.280 632.000 176.400 ;
  LAYER ME1 ;
  RECT 628.460 175.280 632.000 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 619.780 175.280 623.320 176.400 ;
  LAYER ME3 ;
  RECT 619.780 175.280 623.320 176.400 ;
  LAYER ME2 ;
  RECT 619.780 175.280 623.320 176.400 ;
  LAYER ME1 ;
  RECT 619.780 175.280 623.320 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 576.380 175.280 579.920 176.400 ;
  LAYER ME3 ;
  RECT 576.380 175.280 579.920 176.400 ;
  LAYER ME2 ;
  RECT 576.380 175.280 579.920 176.400 ;
  LAYER ME1 ;
  RECT 576.380 175.280 579.920 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 567.700 175.280 571.240 176.400 ;
  LAYER ME3 ;
  RECT 567.700 175.280 571.240 176.400 ;
  LAYER ME2 ;
  RECT 567.700 175.280 571.240 176.400 ;
  LAYER ME1 ;
  RECT 567.700 175.280 571.240 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 559.020 175.280 562.560 176.400 ;
  LAYER ME3 ;
  RECT 559.020 175.280 562.560 176.400 ;
  LAYER ME2 ;
  RECT 559.020 175.280 562.560 176.400 ;
  LAYER ME1 ;
  RECT 559.020 175.280 562.560 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 550.340 175.280 553.880 176.400 ;
  LAYER ME3 ;
  RECT 550.340 175.280 553.880 176.400 ;
  LAYER ME2 ;
  RECT 550.340 175.280 553.880 176.400 ;
  LAYER ME1 ;
  RECT 550.340 175.280 553.880 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 541.660 175.280 545.200 176.400 ;
  LAYER ME3 ;
  RECT 541.660 175.280 545.200 176.400 ;
  LAYER ME2 ;
  RECT 541.660 175.280 545.200 176.400 ;
  LAYER ME1 ;
  RECT 541.660 175.280 545.200 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 532.980 175.280 536.520 176.400 ;
  LAYER ME3 ;
  RECT 532.980 175.280 536.520 176.400 ;
  LAYER ME2 ;
  RECT 532.980 175.280 536.520 176.400 ;
  LAYER ME1 ;
  RECT 532.980 175.280 536.520 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 489.580 175.280 493.120 176.400 ;
  LAYER ME3 ;
  RECT 489.580 175.280 493.120 176.400 ;
  LAYER ME2 ;
  RECT 489.580 175.280 493.120 176.400 ;
  LAYER ME1 ;
  RECT 489.580 175.280 493.120 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 480.900 175.280 484.440 176.400 ;
  LAYER ME3 ;
  RECT 480.900 175.280 484.440 176.400 ;
  LAYER ME2 ;
  RECT 480.900 175.280 484.440 176.400 ;
  LAYER ME1 ;
  RECT 480.900 175.280 484.440 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 472.220 175.280 475.760 176.400 ;
  LAYER ME3 ;
  RECT 472.220 175.280 475.760 176.400 ;
  LAYER ME2 ;
  RECT 472.220 175.280 475.760 176.400 ;
  LAYER ME1 ;
  RECT 472.220 175.280 475.760 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 463.540 175.280 467.080 176.400 ;
  LAYER ME3 ;
  RECT 463.540 175.280 467.080 176.400 ;
  LAYER ME2 ;
  RECT 463.540 175.280 467.080 176.400 ;
  LAYER ME1 ;
  RECT 463.540 175.280 467.080 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 454.860 175.280 458.400 176.400 ;
  LAYER ME3 ;
  RECT 454.860 175.280 458.400 176.400 ;
  LAYER ME2 ;
  RECT 454.860 175.280 458.400 176.400 ;
  LAYER ME1 ;
  RECT 454.860 175.280 458.400 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 446.180 175.280 449.720 176.400 ;
  LAYER ME3 ;
  RECT 446.180 175.280 449.720 176.400 ;
  LAYER ME2 ;
  RECT 446.180 175.280 449.720 176.400 ;
  LAYER ME1 ;
  RECT 446.180 175.280 449.720 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 402.780 175.280 406.320 176.400 ;
  LAYER ME3 ;
  RECT 402.780 175.280 406.320 176.400 ;
  LAYER ME2 ;
  RECT 402.780 175.280 406.320 176.400 ;
  LAYER ME1 ;
  RECT 402.780 175.280 406.320 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 394.100 175.280 397.640 176.400 ;
  LAYER ME3 ;
  RECT 394.100 175.280 397.640 176.400 ;
  LAYER ME2 ;
  RECT 394.100 175.280 397.640 176.400 ;
  LAYER ME1 ;
  RECT 394.100 175.280 397.640 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 385.420 175.280 388.960 176.400 ;
  LAYER ME3 ;
  RECT 385.420 175.280 388.960 176.400 ;
  LAYER ME2 ;
  RECT 385.420 175.280 388.960 176.400 ;
  LAYER ME1 ;
  RECT 385.420 175.280 388.960 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 376.740 175.280 380.280 176.400 ;
  LAYER ME3 ;
  RECT 376.740 175.280 380.280 176.400 ;
  LAYER ME2 ;
  RECT 376.740 175.280 380.280 176.400 ;
  LAYER ME1 ;
  RECT 376.740 175.280 380.280 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 368.060 175.280 371.600 176.400 ;
  LAYER ME3 ;
  RECT 368.060 175.280 371.600 176.400 ;
  LAYER ME2 ;
  RECT 368.060 175.280 371.600 176.400 ;
  LAYER ME1 ;
  RECT 368.060 175.280 371.600 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 359.380 175.280 362.920 176.400 ;
  LAYER ME3 ;
  RECT 359.380 175.280 362.920 176.400 ;
  LAYER ME2 ;
  RECT 359.380 175.280 362.920 176.400 ;
  LAYER ME1 ;
  RECT 359.380 175.280 362.920 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 315.980 175.280 319.520 176.400 ;
  LAYER ME3 ;
  RECT 315.980 175.280 319.520 176.400 ;
  LAYER ME2 ;
  RECT 315.980 175.280 319.520 176.400 ;
  LAYER ME1 ;
  RECT 315.980 175.280 319.520 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 307.300 175.280 310.840 176.400 ;
  LAYER ME3 ;
  RECT 307.300 175.280 310.840 176.400 ;
  LAYER ME2 ;
  RECT 307.300 175.280 310.840 176.400 ;
  LAYER ME1 ;
  RECT 307.300 175.280 310.840 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 298.620 175.280 302.160 176.400 ;
  LAYER ME3 ;
  RECT 298.620 175.280 302.160 176.400 ;
  LAYER ME2 ;
  RECT 298.620 175.280 302.160 176.400 ;
  LAYER ME1 ;
  RECT 298.620 175.280 302.160 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 289.940 175.280 293.480 176.400 ;
  LAYER ME3 ;
  RECT 289.940 175.280 293.480 176.400 ;
  LAYER ME2 ;
  RECT 289.940 175.280 293.480 176.400 ;
  LAYER ME1 ;
  RECT 289.940 175.280 293.480 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 281.260 175.280 284.800 176.400 ;
  LAYER ME3 ;
  RECT 281.260 175.280 284.800 176.400 ;
  LAYER ME2 ;
  RECT 281.260 175.280 284.800 176.400 ;
  LAYER ME1 ;
  RECT 281.260 175.280 284.800 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 272.580 175.280 276.120 176.400 ;
  LAYER ME3 ;
  RECT 272.580 175.280 276.120 176.400 ;
  LAYER ME2 ;
  RECT 272.580 175.280 276.120 176.400 ;
  LAYER ME1 ;
  RECT 272.580 175.280 276.120 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 229.180 175.280 232.720 176.400 ;
  LAYER ME3 ;
  RECT 229.180 175.280 232.720 176.400 ;
  LAYER ME2 ;
  RECT 229.180 175.280 232.720 176.400 ;
  LAYER ME1 ;
  RECT 229.180 175.280 232.720 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 220.500 175.280 224.040 176.400 ;
  LAYER ME3 ;
  RECT 220.500 175.280 224.040 176.400 ;
  LAYER ME2 ;
  RECT 220.500 175.280 224.040 176.400 ;
  LAYER ME1 ;
  RECT 220.500 175.280 224.040 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 211.820 175.280 215.360 176.400 ;
  LAYER ME3 ;
  RECT 211.820 175.280 215.360 176.400 ;
  LAYER ME2 ;
  RECT 211.820 175.280 215.360 176.400 ;
  LAYER ME1 ;
  RECT 211.820 175.280 215.360 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 203.140 175.280 206.680 176.400 ;
  LAYER ME3 ;
  RECT 203.140 175.280 206.680 176.400 ;
  LAYER ME2 ;
  RECT 203.140 175.280 206.680 176.400 ;
  LAYER ME1 ;
  RECT 203.140 175.280 206.680 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 194.460 175.280 198.000 176.400 ;
  LAYER ME3 ;
  RECT 194.460 175.280 198.000 176.400 ;
  LAYER ME2 ;
  RECT 194.460 175.280 198.000 176.400 ;
  LAYER ME1 ;
  RECT 194.460 175.280 198.000 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 185.780 175.280 189.320 176.400 ;
  LAYER ME3 ;
  RECT 185.780 175.280 189.320 176.400 ;
  LAYER ME2 ;
  RECT 185.780 175.280 189.320 176.400 ;
  LAYER ME1 ;
  RECT 185.780 175.280 189.320 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 142.380 175.280 145.920 176.400 ;
  LAYER ME3 ;
  RECT 142.380 175.280 145.920 176.400 ;
  LAYER ME2 ;
  RECT 142.380 175.280 145.920 176.400 ;
  LAYER ME1 ;
  RECT 142.380 175.280 145.920 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 133.700 175.280 137.240 176.400 ;
  LAYER ME3 ;
  RECT 133.700 175.280 137.240 176.400 ;
  LAYER ME2 ;
  RECT 133.700 175.280 137.240 176.400 ;
  LAYER ME1 ;
  RECT 133.700 175.280 137.240 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 125.020 175.280 128.560 176.400 ;
  LAYER ME3 ;
  RECT 125.020 175.280 128.560 176.400 ;
  LAYER ME2 ;
  RECT 125.020 175.280 128.560 176.400 ;
  LAYER ME1 ;
  RECT 125.020 175.280 128.560 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 116.340 175.280 119.880 176.400 ;
  LAYER ME3 ;
  RECT 116.340 175.280 119.880 176.400 ;
  LAYER ME2 ;
  RECT 116.340 175.280 119.880 176.400 ;
  LAYER ME1 ;
  RECT 116.340 175.280 119.880 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 107.660 175.280 111.200 176.400 ;
  LAYER ME3 ;
  RECT 107.660 175.280 111.200 176.400 ;
  LAYER ME2 ;
  RECT 107.660 175.280 111.200 176.400 ;
  LAYER ME1 ;
  RECT 107.660 175.280 111.200 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 98.980 175.280 102.520 176.400 ;
  LAYER ME3 ;
  RECT 98.980 175.280 102.520 176.400 ;
  LAYER ME2 ;
  RECT 98.980 175.280 102.520 176.400 ;
  LAYER ME1 ;
  RECT 98.980 175.280 102.520 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 55.580 175.280 59.120 176.400 ;
  LAYER ME3 ;
  RECT 55.580 175.280 59.120 176.400 ;
  LAYER ME2 ;
  RECT 55.580 175.280 59.120 176.400 ;
  LAYER ME1 ;
  RECT 55.580 175.280 59.120 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 46.900 175.280 50.440 176.400 ;
  LAYER ME3 ;
  RECT 46.900 175.280 50.440 176.400 ;
  LAYER ME2 ;
  RECT 46.900 175.280 50.440 176.400 ;
  LAYER ME1 ;
  RECT 46.900 175.280 50.440 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 38.220 175.280 41.760 176.400 ;
  LAYER ME3 ;
  RECT 38.220 175.280 41.760 176.400 ;
  LAYER ME2 ;
  RECT 38.220 175.280 41.760 176.400 ;
  LAYER ME1 ;
  RECT 38.220 175.280 41.760 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 29.540 175.280 33.080 176.400 ;
  LAYER ME3 ;
  RECT 29.540 175.280 33.080 176.400 ;
  LAYER ME2 ;
  RECT 29.540 175.280 33.080 176.400 ;
  LAYER ME1 ;
  RECT 29.540 175.280 33.080 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 20.860 175.280 24.400 176.400 ;
  LAYER ME3 ;
  RECT 20.860 175.280 24.400 176.400 ;
  LAYER ME2 ;
  RECT 20.860 175.280 24.400 176.400 ;
  LAYER ME1 ;
  RECT 20.860 175.280 24.400 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 12.180 175.280 15.720 176.400 ;
  LAYER ME3 ;
  RECT 12.180 175.280 15.720 176.400 ;
  LAYER ME2 ;
  RECT 12.180 175.280 15.720 176.400 ;
  LAYER ME1 ;
  RECT 12.180 175.280 15.720 176.400 ;
 END
 PORT
  LAYER ME4 ;
  RECT 975.040 0.000 978.580 1.120 ;
  LAYER ME3 ;
  RECT 975.040 0.000 978.580 1.120 ;
  LAYER ME2 ;
  RECT 975.040 0.000 978.580 1.120 ;
  LAYER ME1 ;
  RECT 975.040 0.000 978.580 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 953.340 0.000 956.880 1.120 ;
  LAYER ME3 ;
  RECT 953.340 0.000 956.880 1.120 ;
  LAYER ME2 ;
  RECT 953.340 0.000 956.880 1.120 ;
  LAYER ME1 ;
  RECT 953.340 0.000 956.880 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 931.640 0.000 935.180 1.120 ;
  LAYER ME3 ;
  RECT 931.640 0.000 935.180 1.120 ;
  LAYER ME2 ;
  RECT 931.640 0.000 935.180 1.120 ;
  LAYER ME1 ;
  RECT 931.640 0.000 935.180 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 904.980 0.000 908.520 1.120 ;
  LAYER ME3 ;
  RECT 904.980 0.000 908.520 1.120 ;
  LAYER ME2 ;
  RECT 904.980 0.000 908.520 1.120 ;
  LAYER ME1 ;
  RECT 904.980 0.000 908.520 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 792.140 0.000 795.680 1.120 ;
  LAYER ME3 ;
  RECT 792.140 0.000 795.680 1.120 ;
  LAYER ME2 ;
  RECT 792.140 0.000 795.680 1.120 ;
  LAYER ME1 ;
  RECT 792.140 0.000 795.680 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 775.400 0.000 778.940 1.120 ;
  LAYER ME3 ;
  RECT 775.400 0.000 778.940 1.120 ;
  LAYER ME2 ;
  RECT 775.400 0.000 778.940 1.120 ;
  LAYER ME1 ;
  RECT 775.400 0.000 778.940 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 748.740 0.000 752.280 1.120 ;
  LAYER ME3 ;
  RECT 748.740 0.000 752.280 1.120 ;
  LAYER ME2 ;
  RECT 748.740 0.000 752.280 1.120 ;
  LAYER ME1 ;
  RECT 748.740 0.000 752.280 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 727.040 0.000 730.580 1.120 ;
  LAYER ME3 ;
  RECT 727.040 0.000 730.580 1.120 ;
  LAYER ME2 ;
  RECT 727.040 0.000 730.580 1.120 ;
  LAYER ME1 ;
  RECT 727.040 0.000 730.580 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 705.340 0.000 708.880 1.120 ;
  LAYER ME3 ;
  RECT 705.340 0.000 708.880 1.120 ;
  LAYER ME2 ;
  RECT 705.340 0.000 708.880 1.120 ;
  LAYER ME1 ;
  RECT 705.340 0.000 708.880 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 678.680 0.000 682.220 1.120 ;
  LAYER ME3 ;
  RECT 678.680 0.000 682.220 1.120 ;
  LAYER ME2 ;
  RECT 678.680 0.000 682.220 1.120 ;
  LAYER ME1 ;
  RECT 678.680 0.000 682.220 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 565.840 0.000 569.380 1.120 ;
  LAYER ME3 ;
  RECT 565.840 0.000 569.380 1.120 ;
  LAYER ME2 ;
  RECT 565.840 0.000 569.380 1.120 ;
  LAYER ME1 ;
  RECT 565.840 0.000 569.380 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 549.100 0.000 552.640 1.120 ;
  LAYER ME3 ;
  RECT 549.100 0.000 552.640 1.120 ;
  LAYER ME2 ;
  RECT 549.100 0.000 552.640 1.120 ;
  LAYER ME1 ;
  RECT 549.100 0.000 552.640 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 513.140 0.000 516.680 1.120 ;
  LAYER ME3 ;
  RECT 513.140 0.000 516.680 1.120 ;
  LAYER ME2 ;
  RECT 513.140 0.000 516.680 1.120 ;
  LAYER ME1 ;
  RECT 513.140 0.000 516.680 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 504.460 0.000 508.000 1.120 ;
  LAYER ME3 ;
  RECT 504.460 0.000 508.000 1.120 ;
  LAYER ME2 ;
  RECT 504.460 0.000 508.000 1.120 ;
  LAYER ME1 ;
  RECT 504.460 0.000 508.000 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 482.760 0.000 486.300 1.120 ;
  LAYER ME3 ;
  RECT 482.760 0.000 486.300 1.120 ;
  LAYER ME2 ;
  RECT 482.760 0.000 486.300 1.120 ;
  LAYER ME1 ;
  RECT 482.760 0.000 486.300 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 465.400 0.000 468.940 1.120 ;
  LAYER ME3 ;
  RECT 465.400 0.000 468.940 1.120 ;
  LAYER ME2 ;
  RECT 465.400 0.000 468.940 1.120 ;
  LAYER ME1 ;
  RECT 465.400 0.000 468.940 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 366.200 0.000 369.740 1.120 ;
  LAYER ME3 ;
  RECT 366.200 0.000 369.740 1.120 ;
  LAYER ME2 ;
  RECT 366.200 0.000 369.740 1.120 ;
  LAYER ME1 ;
  RECT 366.200 0.000 369.740 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 339.540 0.000 343.080 1.120 ;
  LAYER ME3 ;
  RECT 339.540 0.000 343.080 1.120 ;
  LAYER ME2 ;
  RECT 339.540 0.000 343.080 1.120 ;
  LAYER ME1 ;
  RECT 339.540 0.000 343.080 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 318.460 0.000 322.000 1.120 ;
  LAYER ME3 ;
  RECT 318.460 0.000 322.000 1.120 ;
  LAYER ME2 ;
  RECT 318.460 0.000 322.000 1.120 ;
  LAYER ME1 ;
  RECT 318.460 0.000 322.000 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 296.760 0.000 300.300 1.120 ;
  LAYER ME3 ;
  RECT 296.760 0.000 300.300 1.120 ;
  LAYER ME2 ;
  RECT 296.760 0.000 300.300 1.120 ;
  LAYER ME1 ;
  RECT 296.760 0.000 300.300 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 270.100 0.000 273.640 1.120 ;
  LAYER ME3 ;
  RECT 270.100 0.000 273.640 1.120 ;
  LAYER ME2 ;
  RECT 270.100 0.000 273.640 1.120 ;
  LAYER ME1 ;
  RECT 270.100 0.000 273.640 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 253.360 0.000 256.900 1.120 ;
  LAYER ME3 ;
  RECT 253.360 0.000 256.900 1.120 ;
  LAYER ME2 ;
  RECT 253.360 0.000 256.900 1.120 ;
  LAYER ME1 ;
  RECT 253.360 0.000 256.900 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 139.900 0.000 143.440 1.120 ;
  LAYER ME3 ;
  RECT 139.900 0.000 143.440 1.120 ;
  LAYER ME2 ;
  RECT 139.900 0.000 143.440 1.120 ;
  LAYER ME1 ;
  RECT 139.900 0.000 143.440 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 113.860 0.000 117.400 1.120 ;
  LAYER ME3 ;
  RECT 113.860 0.000 117.400 1.120 ;
  LAYER ME2 ;
  RECT 113.860 0.000 117.400 1.120 ;
  LAYER ME1 ;
  RECT 113.860 0.000 117.400 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 92.160 0.000 95.700 1.120 ;
  LAYER ME3 ;
  RECT 92.160 0.000 95.700 1.120 ;
  LAYER ME2 ;
  RECT 92.160 0.000 95.700 1.120 ;
  LAYER ME1 ;
  RECT 92.160 0.000 95.700 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 70.460 0.000 74.000 1.120 ;
  LAYER ME3 ;
  RECT 70.460 0.000 74.000 1.120 ;
  LAYER ME2 ;
  RECT 70.460 0.000 74.000 1.120 ;
  LAYER ME1 ;
  RECT 70.460 0.000 74.000 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 43.800 0.000 47.340 1.120 ;
  LAYER ME3 ;
  RECT 43.800 0.000 47.340 1.120 ;
  LAYER ME2 ;
  RECT 43.800 0.000 47.340 1.120 ;
  LAYER ME1 ;
  RECT 43.800 0.000 47.340 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 27.060 0.000 30.600 1.120 ;
  LAYER ME3 ;
  RECT 27.060 0.000 30.600 1.120 ;
  LAYER ME2 ;
  RECT 27.060 0.000 30.600 1.120 ;
  LAYER ME1 ;
  RECT 27.060 0.000 30.600 1.120 ;
 END
END GND
PIN DO63
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 980.900 0.000 982.020 1.120 ;
  LAYER ME3 ;
  RECT 980.900 0.000 982.020 1.120 ;
  LAYER ME2 ;
  RECT 980.900 0.000 982.020 1.120 ;
  LAYER ME1 ;
  RECT 980.900 0.000 982.020 1.120 ;
 END
END DO63
PIN DI63
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 972.840 0.000 973.960 1.120 ;
  LAYER ME3 ;
  RECT 972.840 0.000 973.960 1.120 ;
  LAYER ME2 ;
  RECT 972.840 0.000 973.960 1.120 ;
  LAYER ME1 ;
  RECT 972.840 0.000 973.960 1.120 ;
 END
END DI63
PIN DO62
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 967.880 0.000 969.000 1.120 ;
  LAYER ME3 ;
  RECT 967.880 0.000 969.000 1.120 ;
  LAYER ME2 ;
  RECT 967.880 0.000 969.000 1.120 ;
  LAYER ME1 ;
  RECT 967.880 0.000 969.000 1.120 ;
 END
END DO62
PIN DI62
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 959.200 0.000 960.320 1.120 ;
  LAYER ME3 ;
  RECT 959.200 0.000 960.320 1.120 ;
  LAYER ME2 ;
  RECT 959.200 0.000 960.320 1.120 ;
  LAYER ME1 ;
  RECT 959.200 0.000 960.320 1.120 ;
 END
END DI62
PIN DO61
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 951.140 0.000 952.260 1.120 ;
  LAYER ME3 ;
  RECT 951.140 0.000 952.260 1.120 ;
  LAYER ME2 ;
  RECT 951.140 0.000 952.260 1.120 ;
  LAYER ME1 ;
  RECT 951.140 0.000 952.260 1.120 ;
 END
END DO61
PIN DI61
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 942.460 0.000 943.580 1.120 ;
  LAYER ME3 ;
  RECT 942.460 0.000 943.580 1.120 ;
  LAYER ME2 ;
  RECT 942.460 0.000 943.580 1.120 ;
  LAYER ME1 ;
  RECT 942.460 0.000 943.580 1.120 ;
 END
END DI61
PIN DO60
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 937.500 0.000 938.620 1.120 ;
  LAYER ME3 ;
  RECT 937.500 0.000 938.620 1.120 ;
  LAYER ME2 ;
  RECT 937.500 0.000 938.620 1.120 ;
  LAYER ME1 ;
  RECT 937.500 0.000 938.620 1.120 ;
 END
END DO60
PIN DI60
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 929.440 0.000 930.560 1.120 ;
  LAYER ME3 ;
  RECT 929.440 0.000 930.560 1.120 ;
  LAYER ME2 ;
  RECT 929.440 0.000 930.560 1.120 ;
  LAYER ME1 ;
  RECT 929.440 0.000 930.560 1.120 ;
 END
END DI60
PIN DO59
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 924.480 0.000 925.600 1.120 ;
  LAYER ME3 ;
  RECT 924.480 0.000 925.600 1.120 ;
  LAYER ME2 ;
  RECT 924.480 0.000 925.600 1.120 ;
  LAYER ME1 ;
  RECT 924.480 0.000 925.600 1.120 ;
 END
END DO59
PIN DI59
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 915.800 0.000 916.920 1.120 ;
  LAYER ME3 ;
  RECT 915.800 0.000 916.920 1.120 ;
  LAYER ME2 ;
  RECT 915.800 0.000 916.920 1.120 ;
  LAYER ME1 ;
  RECT 915.800 0.000 916.920 1.120 ;
 END
END DI59
PIN DO58
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 911.460 0.000 912.580 1.120 ;
  LAYER ME3 ;
  RECT 911.460 0.000 912.580 1.120 ;
  LAYER ME2 ;
  RECT 911.460 0.000 912.580 1.120 ;
  LAYER ME1 ;
  RECT 911.460 0.000 912.580 1.120 ;
 END
END DO58
PIN DI58
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 902.780 0.000 903.900 1.120 ;
  LAYER ME3 ;
  RECT 902.780 0.000 903.900 1.120 ;
  LAYER ME2 ;
  RECT 902.780 0.000 903.900 1.120 ;
  LAYER ME1 ;
  RECT 902.780 0.000 903.900 1.120 ;
 END
END DI58
PIN DO57
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 894.720 0.000 895.840 1.120 ;
  LAYER ME3 ;
  RECT 894.720 0.000 895.840 1.120 ;
  LAYER ME2 ;
  RECT 894.720 0.000 895.840 1.120 ;
  LAYER ME1 ;
  RECT 894.720 0.000 895.840 1.120 ;
 END
END DO57
PIN DI57
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 886.040 0.000 887.160 1.120 ;
  LAYER ME3 ;
  RECT 886.040 0.000 887.160 1.120 ;
  LAYER ME2 ;
  RECT 886.040 0.000 887.160 1.120 ;
  LAYER ME1 ;
  RECT 886.040 0.000 887.160 1.120 ;
 END
END DI57
PIN DO56
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 881.080 0.000 882.200 1.120 ;
  LAYER ME3 ;
  RECT 881.080 0.000 882.200 1.120 ;
  LAYER ME2 ;
  RECT 881.080 0.000 882.200 1.120 ;
  LAYER ME1 ;
  RECT 881.080 0.000 882.200 1.120 ;
 END
END DO56
PIN DI56
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 873.020 0.000 874.140 1.120 ;
  LAYER ME3 ;
  RECT 873.020 0.000 874.140 1.120 ;
  LAYER ME2 ;
  RECT 873.020 0.000 874.140 1.120 ;
  LAYER ME1 ;
  RECT 873.020 0.000 874.140 1.120 ;
 END
END DI56
PIN DO55
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 868.060 0.000 869.180 1.120 ;
  LAYER ME3 ;
  RECT 868.060 0.000 869.180 1.120 ;
  LAYER ME2 ;
  RECT 868.060 0.000 869.180 1.120 ;
  LAYER ME1 ;
  RECT 868.060 0.000 869.180 1.120 ;
 END
END DO55
PIN DI55
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 859.380 0.000 860.500 1.120 ;
  LAYER ME3 ;
  RECT 859.380 0.000 860.500 1.120 ;
  LAYER ME2 ;
  RECT 859.380 0.000 860.500 1.120 ;
  LAYER ME1 ;
  RECT 859.380 0.000 860.500 1.120 ;
 END
END DI55
PIN DO54
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 854.420 0.000 855.540 1.120 ;
  LAYER ME3 ;
  RECT 854.420 0.000 855.540 1.120 ;
  LAYER ME2 ;
  RECT 854.420 0.000 855.540 1.120 ;
  LAYER ME1 ;
  RECT 854.420 0.000 855.540 1.120 ;
 END
END DO54
PIN DI54
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 846.360 0.000 847.480 1.120 ;
  LAYER ME3 ;
  RECT 846.360 0.000 847.480 1.120 ;
  LAYER ME2 ;
  RECT 846.360 0.000 847.480 1.120 ;
  LAYER ME1 ;
  RECT 846.360 0.000 847.480 1.120 ;
 END
END DI54
PIN DO53
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 837.680 0.000 838.800 1.120 ;
  LAYER ME3 ;
  RECT 837.680 0.000 838.800 1.120 ;
  LAYER ME2 ;
  RECT 837.680 0.000 838.800 1.120 ;
  LAYER ME1 ;
  RECT 837.680 0.000 838.800 1.120 ;
 END
END DO53
PIN DI53
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 829.620 0.000 830.740 1.120 ;
  LAYER ME3 ;
  RECT 829.620 0.000 830.740 1.120 ;
  LAYER ME2 ;
  RECT 829.620 0.000 830.740 1.120 ;
  LAYER ME1 ;
  RECT 829.620 0.000 830.740 1.120 ;
 END
END DI53
PIN DO52
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 824.660 0.000 825.780 1.120 ;
  LAYER ME3 ;
  RECT 824.660 0.000 825.780 1.120 ;
  LAYER ME2 ;
  RECT 824.660 0.000 825.780 1.120 ;
  LAYER ME1 ;
  RECT 824.660 0.000 825.780 1.120 ;
 END
END DO52
PIN DI52
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 815.980 0.000 817.100 1.120 ;
  LAYER ME3 ;
  RECT 815.980 0.000 817.100 1.120 ;
  LAYER ME2 ;
  RECT 815.980 0.000 817.100 1.120 ;
  LAYER ME1 ;
  RECT 815.980 0.000 817.100 1.120 ;
 END
END DI52
PIN DO51
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 811.640 0.000 812.760 1.120 ;
  LAYER ME3 ;
  RECT 811.640 0.000 812.760 1.120 ;
  LAYER ME2 ;
  RECT 811.640 0.000 812.760 1.120 ;
  LAYER ME1 ;
  RECT 811.640 0.000 812.760 1.120 ;
 END
END DO51
PIN DI51
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 802.960 0.000 804.080 1.120 ;
  LAYER ME3 ;
  RECT 802.960 0.000 804.080 1.120 ;
  LAYER ME2 ;
  RECT 802.960 0.000 804.080 1.120 ;
  LAYER ME1 ;
  RECT 802.960 0.000 804.080 1.120 ;
 END
END DI51
PIN DO50
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 798.000 0.000 799.120 1.120 ;
  LAYER ME3 ;
  RECT 798.000 0.000 799.120 1.120 ;
  LAYER ME2 ;
  RECT 798.000 0.000 799.120 1.120 ;
  LAYER ME1 ;
  RECT 798.000 0.000 799.120 1.120 ;
 END
END DO50
PIN DI50
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 789.940 0.000 791.060 1.120 ;
  LAYER ME3 ;
  RECT 789.940 0.000 791.060 1.120 ;
  LAYER ME2 ;
  RECT 789.940 0.000 791.060 1.120 ;
  LAYER ME1 ;
  RECT 789.940 0.000 791.060 1.120 ;
 END
END DI50
PIN DO49
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 781.260 0.000 782.380 1.120 ;
  LAYER ME3 ;
  RECT 781.260 0.000 782.380 1.120 ;
  LAYER ME2 ;
  RECT 781.260 0.000 782.380 1.120 ;
  LAYER ME1 ;
  RECT 781.260 0.000 782.380 1.120 ;
 END
END DO49
PIN DI49
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 773.200 0.000 774.320 1.120 ;
  LAYER ME3 ;
  RECT 773.200 0.000 774.320 1.120 ;
  LAYER ME2 ;
  RECT 773.200 0.000 774.320 1.120 ;
  LAYER ME1 ;
  RECT 773.200 0.000 774.320 1.120 ;
 END
END DI49
PIN DO48
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 768.240 0.000 769.360 1.120 ;
  LAYER ME3 ;
  RECT 768.240 0.000 769.360 1.120 ;
  LAYER ME2 ;
  RECT 768.240 0.000 769.360 1.120 ;
  LAYER ME1 ;
  RECT 768.240 0.000 769.360 1.120 ;
 END
END DO48
PIN DI48
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 759.560 0.000 760.680 1.120 ;
  LAYER ME3 ;
  RECT 759.560 0.000 760.680 1.120 ;
  LAYER ME2 ;
  RECT 759.560 0.000 760.680 1.120 ;
  LAYER ME1 ;
  RECT 759.560 0.000 760.680 1.120 ;
 END
END DI48
PIN DO47
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 754.600 0.000 755.720 1.120 ;
  LAYER ME3 ;
  RECT 754.600 0.000 755.720 1.120 ;
  LAYER ME2 ;
  RECT 754.600 0.000 755.720 1.120 ;
  LAYER ME1 ;
  RECT 754.600 0.000 755.720 1.120 ;
 END
END DO47
PIN DI47
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 746.540 0.000 747.660 1.120 ;
  LAYER ME3 ;
  RECT 746.540 0.000 747.660 1.120 ;
  LAYER ME2 ;
  RECT 746.540 0.000 747.660 1.120 ;
  LAYER ME1 ;
  RECT 746.540 0.000 747.660 1.120 ;
 END
END DI47
PIN DO46
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 741.580 0.000 742.700 1.120 ;
  LAYER ME3 ;
  RECT 741.580 0.000 742.700 1.120 ;
  LAYER ME2 ;
  RECT 741.580 0.000 742.700 1.120 ;
  LAYER ME1 ;
  RECT 741.580 0.000 742.700 1.120 ;
 END
END DO46
PIN DI46
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 732.900 0.000 734.020 1.120 ;
  LAYER ME3 ;
  RECT 732.900 0.000 734.020 1.120 ;
  LAYER ME2 ;
  RECT 732.900 0.000 734.020 1.120 ;
  LAYER ME1 ;
  RECT 732.900 0.000 734.020 1.120 ;
 END
END DI46
PIN DO45
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 724.840 0.000 725.960 1.120 ;
  LAYER ME3 ;
  RECT 724.840 0.000 725.960 1.120 ;
  LAYER ME2 ;
  RECT 724.840 0.000 725.960 1.120 ;
  LAYER ME1 ;
  RECT 724.840 0.000 725.960 1.120 ;
 END
END DO45
PIN DI45
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 716.780 0.000 717.900 1.120 ;
  LAYER ME3 ;
  RECT 716.780 0.000 717.900 1.120 ;
  LAYER ME2 ;
  RECT 716.780 0.000 717.900 1.120 ;
  LAYER ME1 ;
  RECT 716.780 0.000 717.900 1.120 ;
 END
END DI45
PIN DO44
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 711.820 0.000 712.940 1.120 ;
  LAYER ME3 ;
  RECT 711.820 0.000 712.940 1.120 ;
  LAYER ME2 ;
  RECT 711.820 0.000 712.940 1.120 ;
  LAYER ME1 ;
  RECT 711.820 0.000 712.940 1.120 ;
 END
END DO44
PIN DI44
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 703.140 0.000 704.260 1.120 ;
  LAYER ME3 ;
  RECT 703.140 0.000 704.260 1.120 ;
  LAYER ME2 ;
  RECT 703.140 0.000 704.260 1.120 ;
  LAYER ME1 ;
  RECT 703.140 0.000 704.260 1.120 ;
 END
END DI44
PIN DO43
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 698.180 0.000 699.300 1.120 ;
  LAYER ME3 ;
  RECT 698.180 0.000 699.300 1.120 ;
  LAYER ME2 ;
  RECT 698.180 0.000 699.300 1.120 ;
  LAYER ME1 ;
  RECT 698.180 0.000 699.300 1.120 ;
 END
END DO43
PIN DI43
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 690.120 0.000 691.240 1.120 ;
  LAYER ME3 ;
  RECT 690.120 0.000 691.240 1.120 ;
  LAYER ME2 ;
  RECT 690.120 0.000 691.240 1.120 ;
  LAYER ME1 ;
  RECT 690.120 0.000 691.240 1.120 ;
 END
END DI43
PIN DO42
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 685.160 0.000 686.280 1.120 ;
  LAYER ME3 ;
  RECT 685.160 0.000 686.280 1.120 ;
  LAYER ME2 ;
  RECT 685.160 0.000 686.280 1.120 ;
  LAYER ME1 ;
  RECT 685.160 0.000 686.280 1.120 ;
 END
END DO42
PIN DI42
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 676.480 0.000 677.600 1.120 ;
  LAYER ME3 ;
  RECT 676.480 0.000 677.600 1.120 ;
  LAYER ME2 ;
  RECT 676.480 0.000 677.600 1.120 ;
  LAYER ME1 ;
  RECT 676.480 0.000 677.600 1.120 ;
 END
END DI42
PIN DO41
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 668.420 0.000 669.540 1.120 ;
  LAYER ME3 ;
  RECT 668.420 0.000 669.540 1.120 ;
  LAYER ME2 ;
  RECT 668.420 0.000 669.540 1.120 ;
  LAYER ME1 ;
  RECT 668.420 0.000 669.540 1.120 ;
 END
END DO41
PIN DI41
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 659.740 0.000 660.860 1.120 ;
  LAYER ME3 ;
  RECT 659.740 0.000 660.860 1.120 ;
  LAYER ME2 ;
  RECT 659.740 0.000 660.860 1.120 ;
  LAYER ME1 ;
  RECT 659.740 0.000 660.860 1.120 ;
 END
END DI41
PIN DO40
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 655.400 0.000 656.520 1.120 ;
  LAYER ME3 ;
  RECT 655.400 0.000 656.520 1.120 ;
  LAYER ME2 ;
  RECT 655.400 0.000 656.520 1.120 ;
  LAYER ME1 ;
  RECT 655.400 0.000 656.520 1.120 ;
 END
END DO40
PIN DI40
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 646.720 0.000 647.840 1.120 ;
  LAYER ME3 ;
  RECT 646.720 0.000 647.840 1.120 ;
  LAYER ME2 ;
  RECT 646.720 0.000 647.840 1.120 ;
  LAYER ME1 ;
  RECT 646.720 0.000 647.840 1.120 ;
 END
END DI40
PIN DO39
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 641.760 0.000 642.880 1.120 ;
  LAYER ME3 ;
  RECT 641.760 0.000 642.880 1.120 ;
  LAYER ME2 ;
  RECT 641.760 0.000 642.880 1.120 ;
  LAYER ME1 ;
  RECT 641.760 0.000 642.880 1.120 ;
 END
END DO39
PIN DI39
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 633.700 0.000 634.820 1.120 ;
  LAYER ME3 ;
  RECT 633.700 0.000 634.820 1.120 ;
  LAYER ME2 ;
  RECT 633.700 0.000 634.820 1.120 ;
  LAYER ME1 ;
  RECT 633.700 0.000 634.820 1.120 ;
 END
END DI39
PIN DO38
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 628.740 0.000 629.860 1.120 ;
  LAYER ME3 ;
  RECT 628.740 0.000 629.860 1.120 ;
  LAYER ME2 ;
  RECT 628.740 0.000 629.860 1.120 ;
  LAYER ME1 ;
  RECT 628.740 0.000 629.860 1.120 ;
 END
END DO38
PIN DI38
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 620.060 0.000 621.180 1.120 ;
  LAYER ME3 ;
  RECT 620.060 0.000 621.180 1.120 ;
  LAYER ME2 ;
  RECT 620.060 0.000 621.180 1.120 ;
  LAYER ME1 ;
  RECT 620.060 0.000 621.180 1.120 ;
 END
END DI38
PIN DO37
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 612.000 0.000 613.120 1.120 ;
  LAYER ME3 ;
  RECT 612.000 0.000 613.120 1.120 ;
  LAYER ME2 ;
  RECT 612.000 0.000 613.120 1.120 ;
  LAYER ME1 ;
  RECT 612.000 0.000 613.120 1.120 ;
 END
END DO37
PIN DI37
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 603.320 0.000 604.440 1.120 ;
  LAYER ME3 ;
  RECT 603.320 0.000 604.440 1.120 ;
  LAYER ME2 ;
  RECT 603.320 0.000 604.440 1.120 ;
  LAYER ME1 ;
  RECT 603.320 0.000 604.440 1.120 ;
 END
END DI37
PIN DO36
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 598.360 0.000 599.480 1.120 ;
  LAYER ME3 ;
  RECT 598.360 0.000 599.480 1.120 ;
  LAYER ME2 ;
  RECT 598.360 0.000 599.480 1.120 ;
  LAYER ME1 ;
  RECT 598.360 0.000 599.480 1.120 ;
 END
END DO36
PIN DI36
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 590.300 0.000 591.420 1.120 ;
  LAYER ME3 ;
  RECT 590.300 0.000 591.420 1.120 ;
  LAYER ME2 ;
  RECT 590.300 0.000 591.420 1.120 ;
  LAYER ME1 ;
  RECT 590.300 0.000 591.420 1.120 ;
 END
END DI36
PIN DO35
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 585.340 0.000 586.460 1.120 ;
  LAYER ME3 ;
  RECT 585.340 0.000 586.460 1.120 ;
  LAYER ME2 ;
  RECT 585.340 0.000 586.460 1.120 ;
  LAYER ME1 ;
  RECT 585.340 0.000 586.460 1.120 ;
 END
END DO35
PIN DI35
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 576.660 0.000 577.780 1.120 ;
  LAYER ME3 ;
  RECT 576.660 0.000 577.780 1.120 ;
  LAYER ME2 ;
  RECT 576.660 0.000 577.780 1.120 ;
  LAYER ME1 ;
  RECT 576.660 0.000 577.780 1.120 ;
 END
END DI35
PIN DO34
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 572.320 0.000 573.440 1.120 ;
  LAYER ME3 ;
  RECT 572.320 0.000 573.440 1.120 ;
  LAYER ME2 ;
  RECT 572.320 0.000 573.440 1.120 ;
  LAYER ME1 ;
  RECT 572.320 0.000 573.440 1.120 ;
 END
END DO34
PIN DI34
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 563.640 0.000 564.760 1.120 ;
  LAYER ME3 ;
  RECT 563.640 0.000 564.760 1.120 ;
  LAYER ME2 ;
  RECT 563.640 0.000 564.760 1.120 ;
  LAYER ME1 ;
  RECT 563.640 0.000 564.760 1.120 ;
 END
END DI34
PIN DO33
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 555.580 0.000 556.700 1.120 ;
  LAYER ME3 ;
  RECT 555.580 0.000 556.700 1.120 ;
  LAYER ME2 ;
  RECT 555.580 0.000 556.700 1.120 ;
  LAYER ME1 ;
  RECT 555.580 0.000 556.700 1.120 ;
 END
END DO33
PIN DI33
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 546.900 0.000 548.020 1.120 ;
  LAYER ME3 ;
  RECT 546.900 0.000 548.020 1.120 ;
  LAYER ME2 ;
  RECT 546.900 0.000 548.020 1.120 ;
  LAYER ME1 ;
  RECT 546.900 0.000 548.020 1.120 ;
 END
END DI33
PIN DO32
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 541.940 0.000 543.060 1.120 ;
  LAYER ME3 ;
  RECT 541.940 0.000 543.060 1.120 ;
  LAYER ME2 ;
  RECT 541.940 0.000 543.060 1.120 ;
  LAYER ME1 ;
  RECT 541.940 0.000 543.060 1.120 ;
 END
END DO32
PIN DI32
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 533.880 0.000 535.000 1.120 ;
  LAYER ME3 ;
  RECT 533.880 0.000 535.000 1.120 ;
  LAYER ME2 ;
  RECT 533.880 0.000 535.000 1.120 ;
  LAYER ME1 ;
  RECT 533.880 0.000 535.000 1.120 ;
 END
END DI32
PIN A1
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 528.300 0.000 529.420 1.120 ;
  LAYER ME3 ;
  RECT 528.300 0.000 529.420 1.120 ;
  LAYER ME2 ;
  RECT 528.300 0.000 529.420 1.120 ;
  LAYER ME1 ;
  RECT 528.300 0.000 529.420 1.120 ;
 END
END A1
PIN WEB
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER ME4 ;
  RECT 526.440 0.000 527.560 1.120 ;
  LAYER ME3 ;
  RECT 526.440 0.000 527.560 1.120 ;
  LAYER ME2 ;
  RECT 526.440 0.000 527.560 1.120 ;
  LAYER ME1 ;
  RECT 526.440 0.000 527.560 1.120 ;
 END
END WEB
PIN OE
  DIRECTION INPUT ;
  CAPACITANCE 0.033 ;
 PORT
  LAYER ME4 ;
  RECT 521.480 0.000 522.600 1.120 ;
  LAYER ME3 ;
  RECT 521.480 0.000 522.600 1.120 ;
  LAYER ME2 ;
  RECT 521.480 0.000 522.600 1.120 ;
  LAYER ME1 ;
  RECT 521.480 0.000 522.600 1.120 ;
 END
END OE
PIN CS
  DIRECTION INPUT ;
  CAPACITANCE 0.123 ;
 PORT
  LAYER ME4 ;
  RECT 519.620 0.000 520.740 1.120 ;
  LAYER ME3 ;
  RECT 519.620 0.000 520.740 1.120 ;
  LAYER ME2 ;
  RECT 519.620 0.000 520.740 1.120 ;
  LAYER ME1 ;
  RECT 519.620 0.000 520.740 1.120 ;
 END
END CS
PIN A2
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 497.920 0.000 499.040 1.120 ;
  LAYER ME3 ;
  RECT 497.920 0.000 499.040 1.120 ;
  LAYER ME2 ;
  RECT 497.920 0.000 499.040 1.120 ;
  LAYER ME1 ;
  RECT 497.920 0.000 499.040 1.120 ;
 END
END A2
PIN CK
  DIRECTION INPUT ;
  CAPACITANCE 0.063 ;
 PORT
  LAYER ME4 ;
  RECT 494.820 0.000 495.940 1.120 ;
  LAYER ME3 ;
  RECT 494.820 0.000 495.940 1.120 ;
  LAYER ME2 ;
  RECT 494.820 0.000 495.940 1.120 ;
  LAYER ME1 ;
  RECT 494.820 0.000 495.940 1.120 ;
 END
END CK
PIN A0
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 492.340 0.000 493.460 1.120 ;
  LAYER ME3 ;
  RECT 492.340 0.000 493.460 1.120 ;
  LAYER ME2 ;
  RECT 492.340 0.000 493.460 1.120 ;
  LAYER ME1 ;
  RECT 492.340 0.000 493.460 1.120 ;
 END
END A0
PIN A3
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 488.000 0.000 489.120 1.120 ;
  LAYER ME3 ;
  RECT 488.000 0.000 489.120 1.120 ;
  LAYER ME2 ;
  RECT 488.000 0.000 489.120 1.120 ;
  LAYER ME1 ;
  RECT 488.000 0.000 489.120 1.120 ;
 END
END A3
PIN A4
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 480.560 0.000 481.680 1.120 ;
  LAYER ME3 ;
  RECT 480.560 0.000 481.680 1.120 ;
  LAYER ME2 ;
  RECT 480.560 0.000 481.680 1.120 ;
  LAYER ME1 ;
  RECT 480.560 0.000 481.680 1.120 ;
 END
END A4
PIN A5
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 477.460 0.000 478.580 1.120 ;
  LAYER ME3 ;
  RECT 477.460 0.000 478.580 1.120 ;
  LAYER ME2 ;
  RECT 477.460 0.000 478.580 1.120 ;
  LAYER ME1 ;
  RECT 477.460 0.000 478.580 1.120 ;
 END
END A5
PIN A6
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 470.020 0.000 471.140 1.120 ;
  LAYER ME3 ;
  RECT 470.020 0.000 471.140 1.120 ;
  LAYER ME2 ;
  RECT 470.020 0.000 471.140 1.120 ;
  LAYER ME1 ;
  RECT 470.020 0.000 471.140 1.120 ;
 END
END A6
PIN DO31
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 458.860 0.000 459.980 1.120 ;
  LAYER ME3 ;
  RECT 458.860 0.000 459.980 1.120 ;
  LAYER ME2 ;
  RECT 458.860 0.000 459.980 1.120 ;
  LAYER ME1 ;
  RECT 458.860 0.000 459.980 1.120 ;
 END
END DO31
PIN DI31
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 450.800 0.000 451.920 1.120 ;
  LAYER ME3 ;
  RECT 450.800 0.000 451.920 1.120 ;
  LAYER ME2 ;
  RECT 450.800 0.000 451.920 1.120 ;
  LAYER ME1 ;
  RECT 450.800 0.000 451.920 1.120 ;
 END
END DI31
PIN DO30
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 445.840 0.000 446.960 1.120 ;
  LAYER ME3 ;
  RECT 445.840 0.000 446.960 1.120 ;
  LAYER ME2 ;
  RECT 445.840 0.000 446.960 1.120 ;
  LAYER ME1 ;
  RECT 445.840 0.000 446.960 1.120 ;
 END
END DO30
PIN DI30
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 437.160 0.000 438.280 1.120 ;
  LAYER ME3 ;
  RECT 437.160 0.000 438.280 1.120 ;
  LAYER ME2 ;
  RECT 437.160 0.000 438.280 1.120 ;
  LAYER ME1 ;
  RECT 437.160 0.000 438.280 1.120 ;
 END
END DI30
PIN DO29
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 429.100 0.000 430.220 1.120 ;
  LAYER ME3 ;
  RECT 429.100 0.000 430.220 1.120 ;
  LAYER ME2 ;
  RECT 429.100 0.000 430.220 1.120 ;
  LAYER ME1 ;
  RECT 429.100 0.000 430.220 1.120 ;
 END
END DO29
PIN DI29
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 420.420 0.000 421.540 1.120 ;
  LAYER ME3 ;
  RECT 420.420 0.000 421.540 1.120 ;
  LAYER ME2 ;
  RECT 420.420 0.000 421.540 1.120 ;
  LAYER ME1 ;
  RECT 420.420 0.000 421.540 1.120 ;
 END
END DI29
PIN DO28
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 415.460 0.000 416.580 1.120 ;
  LAYER ME3 ;
  RECT 415.460 0.000 416.580 1.120 ;
  LAYER ME2 ;
  RECT 415.460 0.000 416.580 1.120 ;
  LAYER ME1 ;
  RECT 415.460 0.000 416.580 1.120 ;
 END
END DO28
PIN DI28
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 407.400 0.000 408.520 1.120 ;
  LAYER ME3 ;
  RECT 407.400 0.000 408.520 1.120 ;
  LAYER ME2 ;
  RECT 407.400 0.000 408.520 1.120 ;
  LAYER ME1 ;
  RECT 407.400 0.000 408.520 1.120 ;
 END
END DI28
PIN DO27
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 402.440 0.000 403.560 1.120 ;
  LAYER ME3 ;
  RECT 402.440 0.000 403.560 1.120 ;
  LAYER ME2 ;
  RECT 402.440 0.000 403.560 1.120 ;
  LAYER ME1 ;
  RECT 402.440 0.000 403.560 1.120 ;
 END
END DO27
PIN DI27
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 393.760 0.000 394.880 1.120 ;
  LAYER ME3 ;
  RECT 393.760 0.000 394.880 1.120 ;
  LAYER ME2 ;
  RECT 393.760 0.000 394.880 1.120 ;
  LAYER ME1 ;
  RECT 393.760 0.000 394.880 1.120 ;
 END
END DI27
PIN DO26
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 389.420 0.000 390.540 1.120 ;
  LAYER ME3 ;
  RECT 389.420 0.000 390.540 1.120 ;
  LAYER ME2 ;
  RECT 389.420 0.000 390.540 1.120 ;
  LAYER ME1 ;
  RECT 389.420 0.000 390.540 1.120 ;
 END
END DO26
PIN DI26
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 380.740 0.000 381.860 1.120 ;
  LAYER ME3 ;
  RECT 380.740 0.000 381.860 1.120 ;
  LAYER ME2 ;
  RECT 380.740 0.000 381.860 1.120 ;
  LAYER ME1 ;
  RECT 380.740 0.000 381.860 1.120 ;
 END
END DI26
PIN DO25
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 372.680 0.000 373.800 1.120 ;
  LAYER ME3 ;
  RECT 372.680 0.000 373.800 1.120 ;
  LAYER ME2 ;
  RECT 372.680 0.000 373.800 1.120 ;
  LAYER ME1 ;
  RECT 372.680 0.000 373.800 1.120 ;
 END
END DO25
PIN DI25
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 364.000 0.000 365.120 1.120 ;
  LAYER ME3 ;
  RECT 364.000 0.000 365.120 1.120 ;
  LAYER ME2 ;
  RECT 364.000 0.000 365.120 1.120 ;
  LAYER ME1 ;
  RECT 364.000 0.000 365.120 1.120 ;
 END
END DI25
PIN DO24
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 359.040 0.000 360.160 1.120 ;
  LAYER ME3 ;
  RECT 359.040 0.000 360.160 1.120 ;
  LAYER ME2 ;
  RECT 359.040 0.000 360.160 1.120 ;
  LAYER ME1 ;
  RECT 359.040 0.000 360.160 1.120 ;
 END
END DO24
PIN DI24
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 350.980 0.000 352.100 1.120 ;
  LAYER ME3 ;
  RECT 350.980 0.000 352.100 1.120 ;
  LAYER ME2 ;
  RECT 350.980 0.000 352.100 1.120 ;
  LAYER ME1 ;
  RECT 350.980 0.000 352.100 1.120 ;
 END
END DI24
PIN DO23
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 346.020 0.000 347.140 1.120 ;
  LAYER ME3 ;
  RECT 346.020 0.000 347.140 1.120 ;
  LAYER ME2 ;
  RECT 346.020 0.000 347.140 1.120 ;
  LAYER ME1 ;
  RECT 346.020 0.000 347.140 1.120 ;
 END
END DO23
PIN DI23
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 337.340 0.000 338.460 1.120 ;
  LAYER ME3 ;
  RECT 337.340 0.000 338.460 1.120 ;
  LAYER ME2 ;
  RECT 337.340 0.000 338.460 1.120 ;
  LAYER ME1 ;
  RECT 337.340 0.000 338.460 1.120 ;
 END
END DI23
PIN DO22
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 332.380 0.000 333.500 1.120 ;
  LAYER ME3 ;
  RECT 332.380 0.000 333.500 1.120 ;
  LAYER ME2 ;
  RECT 332.380 0.000 333.500 1.120 ;
  LAYER ME1 ;
  RECT 332.380 0.000 333.500 1.120 ;
 END
END DO22
PIN DI22
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 324.320 0.000 325.440 1.120 ;
  LAYER ME3 ;
  RECT 324.320 0.000 325.440 1.120 ;
  LAYER ME2 ;
  RECT 324.320 0.000 325.440 1.120 ;
  LAYER ME1 ;
  RECT 324.320 0.000 325.440 1.120 ;
 END
END DI22
PIN DO21
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 316.260 0.000 317.380 1.120 ;
  LAYER ME3 ;
  RECT 316.260 0.000 317.380 1.120 ;
  LAYER ME2 ;
  RECT 316.260 0.000 317.380 1.120 ;
  LAYER ME1 ;
  RECT 316.260 0.000 317.380 1.120 ;
 END
END DO21
PIN DI21
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 307.580 0.000 308.700 1.120 ;
  LAYER ME3 ;
  RECT 307.580 0.000 308.700 1.120 ;
  LAYER ME2 ;
  RECT 307.580 0.000 308.700 1.120 ;
  LAYER ME1 ;
  RECT 307.580 0.000 308.700 1.120 ;
 END
END DI21
PIN DO20
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 302.620 0.000 303.740 1.120 ;
  LAYER ME3 ;
  RECT 302.620 0.000 303.740 1.120 ;
  LAYER ME2 ;
  RECT 302.620 0.000 303.740 1.120 ;
  LAYER ME1 ;
  RECT 302.620 0.000 303.740 1.120 ;
 END
END DO20
PIN DI20
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 294.560 0.000 295.680 1.120 ;
  LAYER ME3 ;
  RECT 294.560 0.000 295.680 1.120 ;
  LAYER ME2 ;
  RECT 294.560 0.000 295.680 1.120 ;
  LAYER ME1 ;
  RECT 294.560 0.000 295.680 1.120 ;
 END
END DI20
PIN DO19
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 289.600 0.000 290.720 1.120 ;
  LAYER ME3 ;
  RECT 289.600 0.000 290.720 1.120 ;
  LAYER ME2 ;
  RECT 289.600 0.000 290.720 1.120 ;
  LAYER ME1 ;
  RECT 289.600 0.000 290.720 1.120 ;
 END
END DO19
PIN DI19
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 280.920 0.000 282.040 1.120 ;
  LAYER ME3 ;
  RECT 280.920 0.000 282.040 1.120 ;
  LAYER ME2 ;
  RECT 280.920 0.000 282.040 1.120 ;
  LAYER ME1 ;
  RECT 280.920 0.000 282.040 1.120 ;
 END
END DI19
PIN DO18
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 275.960 0.000 277.080 1.120 ;
  LAYER ME3 ;
  RECT 275.960 0.000 277.080 1.120 ;
  LAYER ME2 ;
  RECT 275.960 0.000 277.080 1.120 ;
  LAYER ME1 ;
  RECT 275.960 0.000 277.080 1.120 ;
 END
END DO18
PIN DI18
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 267.900 0.000 269.020 1.120 ;
  LAYER ME3 ;
  RECT 267.900 0.000 269.020 1.120 ;
  LAYER ME2 ;
  RECT 267.900 0.000 269.020 1.120 ;
  LAYER ME1 ;
  RECT 267.900 0.000 269.020 1.120 ;
 END
END DI18
PIN DO17
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 259.220 0.000 260.340 1.120 ;
  LAYER ME3 ;
  RECT 259.220 0.000 260.340 1.120 ;
  LAYER ME2 ;
  RECT 259.220 0.000 260.340 1.120 ;
  LAYER ME1 ;
  RECT 259.220 0.000 260.340 1.120 ;
 END
END DO17
PIN DI17
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 251.160 0.000 252.280 1.120 ;
  LAYER ME3 ;
  RECT 251.160 0.000 252.280 1.120 ;
  LAYER ME2 ;
  RECT 251.160 0.000 252.280 1.120 ;
  LAYER ME1 ;
  RECT 251.160 0.000 252.280 1.120 ;
 END
END DI17
PIN DO16
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 246.200 0.000 247.320 1.120 ;
  LAYER ME3 ;
  RECT 246.200 0.000 247.320 1.120 ;
  LAYER ME2 ;
  RECT 246.200 0.000 247.320 1.120 ;
  LAYER ME1 ;
  RECT 246.200 0.000 247.320 1.120 ;
 END
END DO16
PIN DI16
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 237.520 0.000 238.640 1.120 ;
  LAYER ME3 ;
  RECT 237.520 0.000 238.640 1.120 ;
  LAYER ME2 ;
  RECT 237.520 0.000 238.640 1.120 ;
  LAYER ME1 ;
  RECT 237.520 0.000 238.640 1.120 ;
 END
END DI16
PIN DO15
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 233.180 0.000 234.300 1.120 ;
  LAYER ME3 ;
  RECT 233.180 0.000 234.300 1.120 ;
  LAYER ME2 ;
  RECT 233.180 0.000 234.300 1.120 ;
  LAYER ME1 ;
  RECT 233.180 0.000 234.300 1.120 ;
 END
END DO15
PIN DI15
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 224.500 0.000 225.620 1.120 ;
  LAYER ME3 ;
  RECT 224.500 0.000 225.620 1.120 ;
  LAYER ME2 ;
  RECT 224.500 0.000 225.620 1.120 ;
  LAYER ME1 ;
  RECT 224.500 0.000 225.620 1.120 ;
 END
END DI15
PIN DO14
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 219.540 0.000 220.660 1.120 ;
  LAYER ME3 ;
  RECT 219.540 0.000 220.660 1.120 ;
  LAYER ME2 ;
  RECT 219.540 0.000 220.660 1.120 ;
  LAYER ME1 ;
  RECT 219.540 0.000 220.660 1.120 ;
 END
END DO14
PIN DI14
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 211.480 0.000 212.600 1.120 ;
  LAYER ME3 ;
  RECT 211.480 0.000 212.600 1.120 ;
  LAYER ME2 ;
  RECT 211.480 0.000 212.600 1.120 ;
  LAYER ME1 ;
  RECT 211.480 0.000 212.600 1.120 ;
 END
END DI14
PIN DO13
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 202.800 0.000 203.920 1.120 ;
  LAYER ME3 ;
  RECT 202.800 0.000 203.920 1.120 ;
  LAYER ME2 ;
  RECT 202.800 0.000 203.920 1.120 ;
  LAYER ME1 ;
  RECT 202.800 0.000 203.920 1.120 ;
 END
END DO13
PIN DI13
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 194.740 0.000 195.860 1.120 ;
  LAYER ME3 ;
  RECT 194.740 0.000 195.860 1.120 ;
  LAYER ME2 ;
  RECT 194.740 0.000 195.860 1.120 ;
  LAYER ME1 ;
  RECT 194.740 0.000 195.860 1.120 ;
 END
END DI13
PIN DO12
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 189.780 0.000 190.900 1.120 ;
  LAYER ME3 ;
  RECT 189.780 0.000 190.900 1.120 ;
  LAYER ME2 ;
  RECT 189.780 0.000 190.900 1.120 ;
  LAYER ME1 ;
  RECT 189.780 0.000 190.900 1.120 ;
 END
END DO12
PIN DI12
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 181.100 0.000 182.220 1.120 ;
  LAYER ME3 ;
  RECT 181.100 0.000 182.220 1.120 ;
  LAYER ME2 ;
  RECT 181.100 0.000 182.220 1.120 ;
  LAYER ME1 ;
  RECT 181.100 0.000 182.220 1.120 ;
 END
END DI12
PIN DO11
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 176.140 0.000 177.260 1.120 ;
  LAYER ME3 ;
  RECT 176.140 0.000 177.260 1.120 ;
  LAYER ME2 ;
  RECT 176.140 0.000 177.260 1.120 ;
  LAYER ME1 ;
  RECT 176.140 0.000 177.260 1.120 ;
 END
END DO11
PIN DI11
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 168.080 0.000 169.200 1.120 ;
  LAYER ME3 ;
  RECT 168.080 0.000 169.200 1.120 ;
  LAYER ME2 ;
  RECT 168.080 0.000 169.200 1.120 ;
  LAYER ME1 ;
  RECT 168.080 0.000 169.200 1.120 ;
 END
END DI11
PIN DO10
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 163.120 0.000 164.240 1.120 ;
  LAYER ME3 ;
  RECT 163.120 0.000 164.240 1.120 ;
  LAYER ME2 ;
  RECT 163.120 0.000 164.240 1.120 ;
  LAYER ME1 ;
  RECT 163.120 0.000 164.240 1.120 ;
 END
END DO10
PIN DI10
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 154.440 0.000 155.560 1.120 ;
  LAYER ME3 ;
  RECT 154.440 0.000 155.560 1.120 ;
  LAYER ME2 ;
  RECT 154.440 0.000 155.560 1.120 ;
  LAYER ME1 ;
  RECT 154.440 0.000 155.560 1.120 ;
 END
END DI10
PIN DO9
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 146.380 0.000 147.500 1.120 ;
  LAYER ME3 ;
  RECT 146.380 0.000 147.500 1.120 ;
  LAYER ME2 ;
  RECT 146.380 0.000 147.500 1.120 ;
  LAYER ME1 ;
  RECT 146.380 0.000 147.500 1.120 ;
 END
END DO9
PIN DI9
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 137.700 0.000 138.820 1.120 ;
  LAYER ME3 ;
  RECT 137.700 0.000 138.820 1.120 ;
  LAYER ME2 ;
  RECT 137.700 0.000 138.820 1.120 ;
  LAYER ME1 ;
  RECT 137.700 0.000 138.820 1.120 ;
 END
END DI9
PIN DO8
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 133.360 0.000 134.480 1.120 ;
  LAYER ME3 ;
  RECT 133.360 0.000 134.480 1.120 ;
  LAYER ME2 ;
  RECT 133.360 0.000 134.480 1.120 ;
  LAYER ME1 ;
  RECT 133.360 0.000 134.480 1.120 ;
 END
END DO8
PIN DI8
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 124.680 0.000 125.800 1.120 ;
  LAYER ME3 ;
  RECT 124.680 0.000 125.800 1.120 ;
  LAYER ME2 ;
  RECT 124.680 0.000 125.800 1.120 ;
  LAYER ME1 ;
  RECT 124.680 0.000 125.800 1.120 ;
 END
END DI8
PIN DO7
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 119.720 0.000 120.840 1.120 ;
  LAYER ME3 ;
  RECT 119.720 0.000 120.840 1.120 ;
  LAYER ME2 ;
  RECT 119.720 0.000 120.840 1.120 ;
  LAYER ME1 ;
  RECT 119.720 0.000 120.840 1.120 ;
 END
END DO7
PIN DI7
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 111.660 0.000 112.780 1.120 ;
  LAYER ME3 ;
  RECT 111.660 0.000 112.780 1.120 ;
  LAYER ME2 ;
  RECT 111.660 0.000 112.780 1.120 ;
  LAYER ME1 ;
  RECT 111.660 0.000 112.780 1.120 ;
 END
END DI7
PIN DO6
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 106.700 0.000 107.820 1.120 ;
  LAYER ME3 ;
  RECT 106.700 0.000 107.820 1.120 ;
  LAYER ME2 ;
  RECT 106.700 0.000 107.820 1.120 ;
  LAYER ME1 ;
  RECT 106.700 0.000 107.820 1.120 ;
 END
END DO6
PIN DI6
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 98.020 0.000 99.140 1.120 ;
  LAYER ME3 ;
  RECT 98.020 0.000 99.140 1.120 ;
  LAYER ME2 ;
  RECT 98.020 0.000 99.140 1.120 ;
  LAYER ME1 ;
  RECT 98.020 0.000 99.140 1.120 ;
 END
END DI6
PIN DO5
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 89.960 0.000 91.080 1.120 ;
  LAYER ME3 ;
  RECT 89.960 0.000 91.080 1.120 ;
  LAYER ME2 ;
  RECT 89.960 0.000 91.080 1.120 ;
  LAYER ME1 ;
  RECT 89.960 0.000 91.080 1.120 ;
 END
END DO5
PIN DI5
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 81.280 0.000 82.400 1.120 ;
  LAYER ME3 ;
  RECT 81.280 0.000 82.400 1.120 ;
  LAYER ME2 ;
  RECT 81.280 0.000 82.400 1.120 ;
  LAYER ME1 ;
  RECT 81.280 0.000 82.400 1.120 ;
 END
END DI5
PIN DO4
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 76.320 0.000 77.440 1.120 ;
  LAYER ME3 ;
  RECT 76.320 0.000 77.440 1.120 ;
  LAYER ME2 ;
  RECT 76.320 0.000 77.440 1.120 ;
  LAYER ME1 ;
  RECT 76.320 0.000 77.440 1.120 ;
 END
END DO4
PIN DI4
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 68.260 0.000 69.380 1.120 ;
  LAYER ME3 ;
  RECT 68.260 0.000 69.380 1.120 ;
  LAYER ME2 ;
  RECT 68.260 0.000 69.380 1.120 ;
  LAYER ME1 ;
  RECT 68.260 0.000 69.380 1.120 ;
 END
END DI4
PIN DO3
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 63.300 0.000 64.420 1.120 ;
  LAYER ME3 ;
  RECT 63.300 0.000 64.420 1.120 ;
  LAYER ME2 ;
  RECT 63.300 0.000 64.420 1.120 ;
  LAYER ME1 ;
  RECT 63.300 0.000 64.420 1.120 ;
 END
END DO3
PIN DI3
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 54.620 0.000 55.740 1.120 ;
  LAYER ME3 ;
  RECT 54.620 0.000 55.740 1.120 ;
  LAYER ME2 ;
  RECT 54.620 0.000 55.740 1.120 ;
  LAYER ME1 ;
  RECT 54.620 0.000 55.740 1.120 ;
 END
END DI3
PIN DO2
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 50.280 0.000 51.400 1.120 ;
  LAYER ME3 ;
  RECT 50.280 0.000 51.400 1.120 ;
  LAYER ME2 ;
  RECT 50.280 0.000 51.400 1.120 ;
  LAYER ME1 ;
  RECT 50.280 0.000 51.400 1.120 ;
 END
END DO2
PIN DI2
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 41.600 0.000 42.720 1.120 ;
  LAYER ME3 ;
  RECT 41.600 0.000 42.720 1.120 ;
  LAYER ME2 ;
  RECT 41.600 0.000 42.720 1.120 ;
  LAYER ME1 ;
  RECT 41.600 0.000 42.720 1.120 ;
 END
END DI2
PIN DO1
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 33.540 0.000 34.660 1.120 ;
  LAYER ME3 ;
  RECT 33.540 0.000 34.660 1.120 ;
  LAYER ME2 ;
  RECT 33.540 0.000 34.660 1.120 ;
  LAYER ME1 ;
  RECT 33.540 0.000 34.660 1.120 ;
 END
END DO1
PIN DI1
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 24.860 0.000 25.980 1.120 ;
  LAYER ME3 ;
  RECT 24.860 0.000 25.980 1.120 ;
  LAYER ME2 ;
  RECT 24.860 0.000 25.980 1.120 ;
  LAYER ME1 ;
  RECT 24.860 0.000 25.980 1.120 ;
 END
END DI1
PIN DO0
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 19.900 0.000 21.020 1.120 ;
  LAYER ME3 ;
  RECT 19.900 0.000 21.020 1.120 ;
  LAYER ME2 ;
  RECT 19.900 0.000 21.020 1.120 ;
  LAYER ME1 ;
  RECT 19.900 0.000 21.020 1.120 ;
 END
END DO0
PIN DI0
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 11.840 0.000 12.960 1.120 ;
  LAYER ME3 ;
  RECT 11.840 0.000 12.960 1.120 ;
  LAYER ME2 ;
  RECT 11.840 0.000 12.960 1.120 ;
  LAYER ME1 ;
  RECT 11.840 0.000 12.960 1.120 ;
 END
END DI0
OBS
  LAYER ME1 SPACING 0.280 ;
  RECT 0.000 0.140 994.480 176.400 ;
  LAYER ME2 SPACING 0.320 ;
  RECT 0.000 0.140 994.480 176.400 ;
  LAYER ME3 SPACING 0.320 ;
  RECT 0.000 0.140 994.480 176.400 ;
  LAYER ME4 SPACING 0.600 ;
  RECT 0.000 0.140 994.480 176.400 ;
  LAYER VI1 ;
  RECT 0.000 0.140 994.480 176.400 ;
  LAYER VI2 ;
  RECT 0.000 0.140 994.480 176.400 ;
  LAYER VI3 ;
  RECT 0.000 0.140 994.480 176.400 ;
END
END Memory_64_128
END LIBRARY



