// ##############################################################
//   You can modify by your own
//   You can modify by your own
//   You can modify by your own
// ##############################################################

module CHIP(
    // input signals
    clk,
    rst_n,
    in_valid, 
    in_valid2,
    
    image,
    template,
    image_size,
	action,
	
    // output signals
    out_valid,
    out_value
);


input            clk, rst_n, in_valid, in_valid2;
input     [7:0]  image;
input     [7:0]  template;
input     [1:0]  image_size;
input     [2:0]  action;

output           out_valid;
output           out_value;

//==================================================================
// reg & wire
//==================================================================
wire             C_clk;
wire             C_rst_n;
wire             C_in_valid;
wire             C_in_valid2;

wire     [7:0]   C_image;
wire     [7:0]   C_template;
wire     [1:0]   C_image_size;
wire     [2:0]   C_action;

wire             C_out_valid;
wire             C_out_value;

//==================================================================
// CORE
//==================================================================
TMIP CORE(
	// input signals
    .clk(C_clk),
    .rst_n(C_rst_n),
    .in_valid(C_in_valid), 
    .in_valid2(C_in_valid2),
    
    .image(C_image),
    .template(C_template),
    .image_size(C_image_size),
	.action(C_action),
	
    // output signals
    .out_valid(C_out_valid),
    .out_value(C_out_value)
);

//==================================================================
// INPUT PAD
// Syntax: XMD PAD_NAME ( .O(CORE_PORT_NAME), .I(CHIP_PORT_NAME), .PU(1'b0), .PD(1'b0), .SMT(1'b0));
//     Ex: XMD    I_CLK ( .O(C_clk),          .I(clk),            .PU(1'b0), .PD(1'b0), .SMT(1'b0));
//==================================================================
// You need to finish this part
XMD I_CLK               ( .O(C_clk),            .I(clk),                .PU(1'b0), .PD(1'b0), .SMT(1'b0));
XMD I_RST               ( .O(C_rst_n),          .I(rst_n),              .PU(1'b0), .PD(1'b0), .SMT(1'b0));
XMD I_IN_VALID          ( .O(C_in_valid),       .I(in_valid),           .PU(1'b0), .PD(1'b0), .SMT(1'b0));
XMD I_IN_VALID2         ( .O(C_in_valid2),      .I(in_valid2),          .PU(1'b0), .PD(1'b0), .SMT(1'b0));
XMD I_IMAGE0            ( .O(C_image[0]),       .I(image[0]),           .PU(1'b0), .PD(1'b0), .SMT(1'b0));
XMD I_IMAGE1            ( .O(C_image[1]),       .I(image[1]),           .PU(1'b0), .PD(1'b0), .SMT(1'b0));
XMD I_IMAGE2            ( .O(C_image[2]),       .I(image[2]),           .PU(1'b0), .PD(1'b0), .SMT(1'b0));
XMD I_IMAGE3            ( .O(C_image[3]),       .I(image[3]),           .PU(1'b0), .PD(1'b0), .SMT(1'b0));
XMD I_IMAGE4            ( .O(C_image[4]),       .I(image[4]),           .PU(1'b0), .PD(1'b0), .SMT(1'b0));
XMD I_IMAGE5            ( .O(C_image[5]),       .I(image[5]),           .PU(1'b0), .PD(1'b0), .SMT(1'b0));
XMD I_IMAGE6            ( .O(C_image[6]),       .I(image[6]),           .PU(1'b0), .PD(1'b0), .SMT(1'b0));
XMD I_IMAGE7            ( .O(C_image[7]),       .I(image[7]),           .PU(1'b0), .PD(1'b0), .SMT(1'b0));

XMD I_TEMPLATE0            ( .O(C_template[0]),       .I(template[0]),           .PU(1'b0), .PD(1'b0), .SMT(1'b0));
XMD I_TEMPLATE1            ( .O(C_template[1]),       .I(template[1]),           .PU(1'b0), .PD(1'b0), .SMT(1'b0));
XMD I_TEMPLATE2            ( .O(C_template[2]),       .I(template[2]),           .PU(1'b0), .PD(1'b0), .SMT(1'b0));
XMD I_TEMPLATE3            ( .O(C_template[3]),       .I(template[3]),           .PU(1'b0), .PD(1'b0), .SMT(1'b0));
XMD I_TEMPLATE4            ( .O(C_template[4]),       .I(template[4]),           .PU(1'b0), .PD(1'b0), .SMT(1'b0));
XMD I_TEMPLATE5            ( .O(C_template[5]),       .I(template[5]),           .PU(1'b0), .PD(1'b0), .SMT(1'b0));
XMD I_TEMPLATE6            ( .O(C_template[6]),       .I(template[6]),           .PU(1'b0), .PD(1'b0), .SMT(1'b0));
XMD I_TEMPLATE7            ( .O(C_template[7]),       .I(template[7]),           .PU(1'b0), .PD(1'b0), .SMT(1'b0));

XMD I_IMG_SIZE0            ( .O(C_image_size[0]),       .I(image_size[0]),           .PU(1'b0), .PD(1'b0), .SMT(1'b0));
XMD I_IMG_SIZE1            ( .O(C_image_size[1]),       .I(image_size[1]),           .PU(1'b0), .PD(1'b0), .SMT(1'b0));

XMD I_ACTION0            ( .O(C_action[0]),       .I(action[0]),           .PU(1'b0), .PD(1'b0), .SMT(1'b0));
XMD I_ACTION1            ( .O(C_action[1]),       .I(action[1]),           .PU(1'b0), .PD(1'b0), .SMT(1'b0));
XMD I_ACTION2            ( .O(C_action[2]),       .I(action[2]),           .PU(1'b0), .PD(1'b0), .SMT(1'b0));
// 25 input
//==================================================================
// OUTPUT PAD
// Syntax: YA2GSD PAD_NAME (.I(CORE_PIN_NAME), .O(PAD_PIN_NAME), .E(1'b1), .E2(1'b1), .E4(1'b1), .E8(1'b0), .SR(1'b0));
//     Ex: YA2GSD  O_VALID (.I(C_out_valid),   .O(out_valid),    .E(1'b1), .E2(1'b1), .E4(1'b1), .E8(1'b0), .SR(1'b0));
//==================================================================
// You need to finish this part
YA2GSD  O_VALID (.I(C_out_valid),   .O(out_valid),    .E(1'b1), .E2(1'b1), .E4(1'b1), .E8(1'b0), .SR(1'b0));
YA2GSD  O_VALUE (.I(C_out_value),   .O(out_value),    .E(1'b1), .E2(1'b1), .E4(1'b1), .E8(1'b0), .SR(1'b0));
// 2 output
//==================================================================
// I/O power 3.3V pads x? (DVDD + DGND)
// Syntax: VCC3IOD/GNDIOD PAD_NAME ();
//    Ex1: VCC3IOD        VDDP0 ();
//    Ex2: GNDIOD         GNDP0 ();
//==================================================================
// You need to finish this part
VCC3IOD        VDDP0 ();
GNDIOD         GNDP0 ();
VCC3IOD        VDDP1 ();
GNDIOD         GNDP1 ();
VCC3IOD        VDDP2 ();
GNDIOD         GNDP2 ();
VCC3IOD        VDDP3 ();
GNDIOD         GNDP3 ();
VCC3IOD        VDDP4 ();
GNDIOD         GNDP4 ();

//==================================================================
// Core power 1.8V pads x? (VDD + GND)
// Syntax: VCCKD/GNDKD PAD_NAME ();
//    Ex1: VCCKD       VDDC0 ();
//    Ex2: GNDKD       GNDC0 ();
//==================================================================
// You need to finish this part
VCCKD VDDC0 ();
GNDKD GNDC0 ();
VCCKD VDDC1 ();
GNDKD GNDC1 ();
VCCKD VDDC2 ();
GNDKD GNDC2 ();
VCCKD VDDC3 ();
GNDKD GNDC3 ();
VCCKD VDDC4 ();
GNDKD GNDC4 ();
endmodule

/////////////////////////////////////////////////////////////
// Created by: Synopsys DC Ultra(TM) in wire load mode
// Version   : T-2022.03
// Date      : Thu Nov 28 12:58:24 2024
/////////////////////////////////////////////////////////////


module TMIP ( clk, rst_n, in_valid, in_valid2, image, template, image_size, 
        action, out_valid, out_value );
  input [7:0] image;
  input [7:0] template;
  input [1:0] image_size;
  input [2:0] action;
  input clk, rst_n, in_valid, in_valid2;
  output out_valid, out_value;
  wire   act_delay2, N1330, act_delay1, N25777, N25778, N25894, PE_N143,
         PE_N142, PE_N141, PE_N140, PE_N139, PE_N138, PE_N137, PE_N136,
         PE_N135, PE_N134, PE_N133, PE_N132, PE_N131, PE_N130, PE_N129,
         PE_N128, PE_N127, PE_N126, PE_N125, PE_N124, PE_N123, PE_N122,
         PE_N121, PE_N120, PE_N119, PE_N118, PE_N117, PE_N116, PE_N115,
         PE_N114, PE_N113, PE_N112, PE_N111, PE_N110, PE_N109, PE_N108,
         PE_N107, PE_N106, PE_N105, PE_N104, PE_N103, PE_N102, PE_N101,
         PE_N100, PE_N99, PE_N98, PE_N97, PE_N96, PE_N95, PE_N94, PE_N93,
         PE_N92, PE_N91, PE_N90, PE_N89, PE_N88, PE_N87, PE_N86, PE_N85,
         PE_N84, PE_N83, PE_N82, PE_N81, PE_N80, PE_N79, PE_N78, PE_N77,
         PE_N76, PE_N75, PE_N74, PE_N73, PE_N72, PE_N71, PE_N70, PE_N69,
         PE_N68, PE_N67, PE_N66, PE_N65, PE_N64, PE_N63, PE_N62, PE_N61,
         PE_N60, PE_N59, PE_N58, PE_N57, PE_N56, PE_N55, PE_N54, PE_N53,
         PE_N52, PE_N51, PE_N50, PE_N49, PE_N48, PE_N47, PE_N46, PE_N45,
         PE_N44, PE_N43, PE_N42, PE_N41, PE_N40, PE_N39, PE_N38, PE_N37,
         PE_N36, PE_N35, PE_N34, PE_N33, PE_N32, PE_N31, PE_N30, PE_N29,
         PE_N28, PE_N27, PE_N26, PE_N25, PE_N24, PE_N23, PE_N22, PE_N21,
         PE_N20, PE_N19, PE_N18, PE_N17, PE_N16, PE_N15, PE_N14, PE_N13,
         PE_N12, PE_N11, PE_N10, PE_N9, PE_N8, PE_N7, PE_N6, PE_N5, PE_N4,
         PE_N3, PE_N2, PE_N1, PE_N0, n11201, n11202, n11203, n11204, n11205,
         n11206, n11207, n11208, n11209, n11210, n11211, n11212, n11213,
         n11214, n11215, n11216, n11217, n11218, n11219, n11220, n11221,
         n11222, n11223, n11224, n11225, n11226, n11227, n11228, n11229,
         n11230, n11231, n11232, n11233, n11234, n11235, n11236, n11237,
         n11238, n11239, n11240, n11241, n11242, n11243, n11244, n11245,
         n11246, n11247, n11248, n11249, n11250, n11251, n11252, n11253,
         n11254, n11255, n11256, n11257, n11258, n11259, n11260, n11261,
         n11262, n11263, n11264, n11265, n11266, n11267, n11268, n11269,
         n11270, n11271, n11272, n11273, n11274, n11275, n11276, n11277,
         n11278, n11279, n11280, n11281, n11282, n11283, n11284, n11285,
         n11286, n11287, n11288, n11289, n11290, n11291, n11292, n11293,
         n11294, n11295, n11296, n11297, n11298, n11299, n11300, n11301,
         n11302, n11303, n11304, n11305, n11306, n11307, n11308, n11309,
         n11310, n11311, n11312, n11313, n11314, n11315, n11316, n11317,
         n11318, n11319, n11320, n11321, n11322, n11323, n11324, n11325,
         n11326, n11327, n11328, n11329, n11330, n11331, n11332, n11333,
         n11334, n11335, n11336, n11337, n11338, n11339, n11340, n11341,
         n11342, n11343, n11344, n11345, n11346, n11347, n11348, n11349,
         n11350, n11351, n11352, n11353, n11354, n11355, n11356, n11357,
         n11358, n11359, n11360, n11361, n11362, n11363, n11364, n11365,
         n11366, n11367, n11368, n11369, n11370, n11371, n11372, n11373,
         n11374, n11375, n11376, n11377, n11378, n11379, n11380, n11381,
         n11382, n11383, n11384, n11385, n11386, n11387, n11388, n11389,
         n11390, n11391, n11392, n11393, n11394, n11395, n11396, n11397,
         n11398, n11399, n11400, n11401, n11402, n11403, n11404, n11405,
         n11406, n11407, n11408, n11409, n11410, n11411, n11412, n11413,
         n11414, n11415, n11416, n11417, n11418, n11419, n11420, n11421,
         n11422, n11423, n11424, n11425, n11426, n11427, n11428, n11429,
         n11430, n11431, n11432, n11433, n11434, n11435, n11436, n11437,
         n11438, n11439, n11440, n11441, n11442, n11443, n11444, n11445,
         n11446, n11447, n11448, n11449, n11450, n11451, n11452, n11453,
         n11454, n11455, n11456, n11457, n11458, n11459, n11460, n11461,
         n11462, n11463, n11464, n11465, n11466, n11467, n11468, n11469,
         n11470, n11471, n11472, n11473, n11474, n11475, n11476, n11477,
         n11478, n11479, n11480, n11481, n11482, n11483, n11484, n11485,
         n11486, n11487, n11488, n11489, n11490, n11491, n11492, n11493,
         n11494, n11495, n11496, n11497, n11498, n11499, n11500, n11501,
         n11502, n11503, n11504, n11505, n11506, n11507, n11508, n11509,
         n11510, n11511, n11512, n11513, n11514, n11515, n11516, n11517,
         n11518, n11519, n11520, n11521, n11522, n11523, n11524, n11525,
         n11526, n11527, n11528, n11529, n11530, n11531, n11532, n11533,
         n11534, n11535, n11536, n11537, n11538, n11539, n11540, n11541,
         n11542, n11543, n11544, n11545, n11546, n11547, n11548, n11549,
         n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11557,
         n11558, n11559, n11560, n11561, n11562, n11563, n11564, n11565,
         n11566, n11567, n11568, n11569, n11570, n11571, n11572, n11573,
         n11574, n11575, n11576, n11577, n11578, n11579, n11580, n11581,
         n11582, n11583, n11584, n11585, n11586, n11587, n11588, n11589,
         n11590, n11591, n11592, n11593, n11594, n11595, n11596, n11597,
         n11598, n11599, n11600, n11601, n11602, n11603, n11604, n11605,
         n11606, n11607, n11608, n11609, n11610, n11611, n11612, n11613,
         n11614, n11615, n11616, n11617, n11618, n11619, n11620, n11621,
         n11622, n11623, n11624, n11625, n11626, n11627, n11628, n11629,
         n11630, n11631, n11632, n11633, n11634, n11635, n11636, n11637,
         n11638, n11639, n11640, n11641, n11642, n11643, n11644, n11645,
         n11646, n11647, n11648, n11649, n11650, n11651, n11652, n11653,
         n11654, n11655, n11656, n11657, n11658, n11659, n11660, n11661,
         n11662, n11663, n11664, n11665, n11666, n11667, n11668, n11669,
         n11670, n11671, n11672, n11673, n11674, n11675, n11676, n11677,
         n11678, n11679, n11680, n11681, n11682, n11683, n11684, n11685,
         n11686, n11687, n11688, n11689, n11690, n11691, n11692, n11693,
         n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701,
         n11702, n11703, n11704, n11705, n11706, n11707, n11708, n11709,
         n11710, n11711, n11712, n11713, n11714, n11715, n11716, n11717,
         n11718, n11719, n11720, n11721, n11722, n11723, n11724, n11725,
         n11726, n11727, n11728, n11729, n11730, n11731, n11732, n11733,
         n11734, n11735, n11736, n11737, n11738, n11739, n11740, n11741,
         n11742, n11743, n11744, n11745, n11746, n11747, n11748, n11749,
         n11750, n11751, n11752, n11753, n11754, n11755, n11756, n11757,
         n11758, n11759, n11760, n11761, n11762, n11763, n11764, n11765,
         n11766, n11767, n11768, n11769, n11770, n11771, n11772, n11773,
         n11774, n11775, n11776, n11777, n11778, n11779, n11780, n11781,
         n11782, n11783, n11784, n11785, n11786, n11787, n11788, n11789,
         n11790, n11791, n11792, n11793, n11794, n11795, n11796, n11797,
         n11798, n11799, n11800, n11801, n11802, n11803, n11804, n11805,
         n11806, n11807, n11808, n11809, n11810, n11811, n11812, n11813,
         n11814, n11815, n11816, n11817, n11818, n11819, n11820, n11821,
         n11822, n11823, n11824, n11825, n11826, n11827, n11828, n11829,
         n11830, n11831, n11832, n11833, n11834, n11835, n11836, n11837,
         n11838, n11839, n11840, n11841, n11842, n11843, n11844, n11845,
         n11846, n11847, n11848, n11849, n11850, n11851, n11852, n11853,
         n11854, n11855, n11856, n11857, n11858, n11859, n11860, n11861,
         n11862, n11863, n11864, n11865, n11866, n11867, n11868, n11869,
         n11870, n11871, n11872, n11873, n11874, n11875, n11876, n11877,
         n11878, n11879, n11880, n11881, n11882, n11883, n11884, n11885,
         n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893,
         n11894, n11895, n11896, n11897, n11898, n11899, n11900, n11901,
         n11902, n11903, n11904, n11905, n11906, n11907, n11908, n11909,
         n11910, n11911, n11912, n11913, n11914, n11915, n11916, n11917,
         n11918, n11919, n11920, n11921, n11922, n11923, n11924, n11925,
         n11926, n11927, n11928, n11929, n11930, n11931, n11932, n11933,
         n11934, n11935, n11936, n11937, n11938, n11939, n11940, n11941,
         n11942, n11943, n11944, n11945, n11946, n11947, n11948, n11949,
         n11950, n11951, n11952, n11953, n11954, n11955, n11956, n11957,
         n11958, n11959, n11960, n11961, n11962, n11963, n11964, n11965,
         n11966, n11967, n11968, n11969, n11970, n11971, n11972, n11973,
         n11974, n11975, n11976, n11977, n11978, n11979, n11980, n11981,
         n11982, n11983, n11984, n11985, n11986, n11987, n11988, n11989,
         n11990, n11991, n11992, n11993, n11994, n11995, n11996, n11997,
         n11998, n11999, n12000, n12001, n12002, n12003, n12004, n12005,
         n12006, n12007, n12008, n12009, n12010, n12011, n12012, n12013,
         n12014, n12015, n12016, n12017, n12018, n12019, n12020, n12021,
         n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029,
         n12030, n12031, n12032, n12033, n12034, n12035, n12036, n12037,
         n12038, n12039, n12040, n12041, n12042, n12043, n12044, n12045,
         n12046, n12047, n12048, n12049, n12050, n12051, n12052, n12053,
         n12054, n12055, n12056, n12057, n12058, n12059, n12060, n12061,
         n12062, n12063, n12064, n12065, n12066, n12067, n12068, n12069,
         n12070, n12071, n12072, n12073, n12074, n12075, n12076, n12077,
         n12078, n12079, n12080, n12081, n12082, n12083, n12084, n12085,
         n12086, n12087, n12088, n12089, n12090, n12091, n12092, n12093,
         n12094, n12095, n12096, n12097, n12098, n12099, n12100, n12101,
         n12102, n12103, n12104, n12105, n12106, n12107, n12108, n12109,
         n12110, n12111, n12112, n12113, n12114, n12115, n12116, n12117,
         n12118, n12119, n12120, n12121, n12122, n12123, n12124, n12125,
         n12126, n12127, n12128, n12129, n12130, n12131, n12132, n12133,
         n12134, n12135, n12136, n12137, n12138, n12139, n12140, n12141,
         n12142, n12143, n12144, n12145, n12146, n12147, n12148, n12149,
         n12150, n12151, n12152, n12153, n12154, n12155, n12156, n12157,
         n12158, n12159, n12160, n12161, n12162, n12163, n12164, n12165,
         n12166, n12167, n12168, n12169, n12170, n12171, n12172, n12173,
         n12174, n12175, n12176, n12177, n12178, n12179, n12180, n12181,
         n12182, n12183, n12184, n12185, n12186, n12187, n12188, n12189,
         n12190, n12191, n12192, n12193, n12194, n12195, n12196, n12197,
         n12198, n12199, n12200, n12201, n12202, n12203, n12204, n12205,
         n12206, n12207, n12208, n12209, n12210, n12211, n12212, n12213,
         n12214, n12215, n12216, n12217, n12218, n12219, n12220, n12221,
         n12222, n12223, n12224, n12225, n12226, n12227, n12228, n12229,
         n12230, n12231, n12232, n12233, n12234, n12235, n12236, n12237,
         n12238, n12239, n12240, n12241, n12242, n12243, n12244, n12245,
         n12246, n12247, n12248, n12249, n12250, n12251, n12252, n12253,
         n12254, n12255, n12256, n12257, n12258, n12259, n12260, n12261,
         n12262, n12263, n12264, n12265, n12266, n12267, n12268, n12269,
         n12270, n12271, n12272, n12273, n12274, n12275, n12276, n12277,
         n12278, n12279, n12280, n12281, n12282, n12283, n12284, n12285,
         n12286, n12287, n12288, n12289, n12290, n12291, n12292, n12293,
         n12294, n12295, n12296, n12297, n12298, n12299, n12300, n12301,
         n12302, n12303, n12304, n12305, n12306, n12307, n12308, n12309,
         n12310, n12311, n12312, n12313, n12314, n12315, n12316, n12317,
         n12318, n12319, n12320, n12321, n12322, n12323, n12324, n12325,
         n12326, n12327, n12328, n12329, n12330, n12331, n12332, n12333,
         n12334, n12335, n12336, n12337, n12338, n12339, n12340, n12341,
         n12342, n12343, n12344, n12345, n12346, n12347, n12348, n12349,
         n12350, n12351, n12352, n12353, n12354, n12355, n12356, n12357,
         n12358, n12359, n12360, n12361, n12362, n12363, n12364, n12365,
         n12366, n12367, n12368, n12369, n12370, n12371, n12372, n12373,
         n12374, n12375, n12376, n12377, n12378, n12379, n12380, n12381,
         n12382, n12383, n12384, n12385, n12386, n12387, n12388, n12389,
         n12390, n12391, n12392, n12393, n12394, n12395, n12396, n12397,
         n12398, n12399, n12400, n12401, n12402, n12403, n12404, n12405,
         n12406, n12407, n12408, n12409, n12410, n12411, n12412, n12413,
         n12414, n12415, n12416, n12417, n12418, n12419, n12420, n12421,
         n12422, n12423, n12424, n12425, n12426, n12427, n12428, n12429,
         n12430, n12431, n12432, n12433, n12434, n12435, n12436, n12437,
         n12438, n12439, n12440, n12441, n12442, n12443, n12444, n12445,
         n12446, n12447, n12448, n12449, n12450, n12451, n12452, n12453,
         n12454, n12455, n12456, n12457, n12458, n12459, n12460, n12461,
         n12462, n12463, n12464, n12465, n12466, n12467, n12468, n12469,
         n12470, n12471, n12472, n12473, n12474, n12475, n12476, n12477,
         n12478, n12479, n12480, n12481, n12482, n12483, n12484, n12485,
         n12486, n12487, n12488, n12489, n12490, n12491, n12492, n12493,
         n12494, n12495, n12496, n12497, n12498, n12499, n12500, n12501,
         n12502, n12503, n12504, n12505, n12506, n12507, n12508, n12509,
         n12510, n12511, n12512, n12513, n12514, n12515, n12516, n12517,
         n12518, n12519, n12520, n12521, n12522, n12523, n12524, n12525,
         n12526, n12527, n12528, n12529, n12530, n12531, n12532, n12533,
         n12534, n12535, n12536, n12537, n12538, n12539, n12540, n12541,
         n12542, n12543, n12544, n12545, n12546, n12547, n12548, n12549,
         n12550, n12551, n12552, n12553, n12554, n12555, n12556, n12557,
         n12558, n12559, n12560, n12561, n12562, n12563, n12564, n12565,
         n12566, n12567, n12568, n12569, n12570, n12571, n12572, n12573,
         n12574, n12575, n12576, n12577, n12578, n12579, n12580, n12581,
         n12582, n12583, n12584, n12585, n12586, n12587, n12588, n12589,
         n12590, n12591, n12592, n12593, n12594, n12595, n12596, n12597,
         n12598, n12599, n12600, n12601, n12602, n12603, n12604, n12605,
         n12606, n12607, n12608, n12609, n12610, n12611, n12612, n12613,
         n12614, n12615, n12616, n12617, n12618, n12619, n12620, n12621,
         n12622, n12623, n12624, n12625, n12626, n12627, n12628, n12629,
         n12630, n12631, n12632, n12633, n12634, n12635, n12636, n12637,
         n12638, n12639, n12640, n12641, n12642, n12643, n12644, n12645,
         n12646, n12647, n12648, n12649, n12650, n12651, n12652, n12653,
         n12654, n12655, n12656, n12657, n12658, n12659, n12660, n12661,
         n12662, n12663, n12664, n12665, n12666, n12667, n12668, n12669,
         n12670, n12671, n12672, n12673, n12674, n12675, n12676, n12677,
         n12678, n12679, n12680, n12681, n12682, n12683, n12684, n12685,
         n12686, n12687, n12688, n12689, n12690, n12691, n12692, n12693,
         n12694, n12695, n12696, n12697, n12698, n12699, n12700, n12701,
         n12702, n12703, n12704, n12705, n12706, n12707, n12708, n12709,
         n12710, n12711, n12712, n12713, n12714, n12715, n12716, n12717,
         n12718, n12719, n12720, n12721, n12722, n12723, n12724, n12725,
         n12726, n12727, n12728, n12729, n12730, n12731, n12732, n12733,
         n12734, n12735, n12736, n12737, n12738, n12739, n12740, n12741,
         n12742, n12743, n12744, n12745, n12746, n12747, n12748, n12749,
         n12750, n12751, n12752, n12753, n12754, n12755, n12756, n12757,
         n12758, n12759, n12760, n12761, n12762, n12763, n12764, n12765,
         n12766, n12767, n12768, n12769, n12770, n12771, n12772, n12773,
         n12774, n12775, n12776, n12777, n12778, n12779, n12780, n12781,
         n12782, n12783, n12784, n12785, n12786, n12787, n12788, n12789,
         n12790, n12791, n12792, n12793, n12794, n12795, n12796, n12797,
         n12798, n12799, n12800, n12801, n12802, n12803, n12804, n12805,
         n12806, n12807, n12808, n12809, n12810, n12811, n12812, n12813,
         n12814, n12815, n12816, n12817, n12818, n12819, n12820, n12821,
         n12822, n12823, n12824, n12825, n12826, n12827, n12828, n12829,
         n12830, n12831, n12832, n12833, n12834, n12835, n12836, n12837,
         n12838, n12839, n12840, n12841, n12842, n12843, n12844, n12845,
         n12846, n12847, n12848, n12849, n12850, n12851, n12852, n12853,
         n12854, n12855, n12856, n12857, n12858, n12859, n12860, n12861,
         n12862, n12863, n12864, n12865, n12866, n12867, n12868, n12869,
         n12870, n12871, n12872, n12873, n12874, n12875, n12876, n12877,
         n12878, n12879, n12880, n12881, n12882, n12883, n12884, n12885,
         n12886, n12887, n12888, n12889, n12890, n12891, n12892, n12893,
         n12894, n12895, n12896, n12897, n12898, n12899, n12900, n12901,
         n12902, n12903, n12904, n12905, n12906, n12907, n12908, n12909,
         n12910, n12911, n12912, n12913, n12914, n12915, n12916, n12917,
         n12918, n12919, n12920, n12921, n12922, n12923, n12924, n12925,
         n12926, n12927, n12928, n12929, n12930, n12931, n12932, n12933,
         n12934, n12935, n12936, n12937, n12938, n12939, n12940, n12941,
         n12942, n12943, n12944, n12945, n12946, n12947, n12948, n12949,
         n12950, n12951, n12952, n12953, n12954, n12955, n12956, n12957,
         n12958, n12959, n12960, n12961, n12962, n12963, n12964, n12965,
         n12966, n12967, n12968, n12969, n12970, n12971, n12972, n12973,
         n12974, n12975, n12976, n12977, n12978, n12979, n12980, n12981,
         n12982, n12983, n12984, n12985, n12986, n12987, n12988, n12989,
         n12990, n12991, n12992, n12993, n12994, n12995, n12996, n12997,
         n12998, n12999, n13000, n13001, n13002, n13003, n13004, n13005,
         n13006, n13007, n13008, n13009, n13010, n13011, n13012, n13013,
         n13014, n13015, n13016, n13017, n13018, n13019, n13020, n13021,
         n13022, n13023, n13024, n13025, n13026, n13027, n13028, n13029,
         n13030, n13031, n13032, n13033, n13034, n13035, n13036, n13037,
         n13038, n13039, n13040, n13041, n13042, n13043, n13044, n13045,
         n13046, n13047, n13048, n13049, n13050, n13051, n13052, n13053,
         n13054, n13055, n13056, n13057, n13058, n13059, n13060, n13061,
         n13062, n13063, n13064, n13065, n13066, n13067, n13068, n13069,
         n13070, n13071, n13072, n13073, n13074, n13075, n13076, n13077,
         n13078, n13079, n13080, n13081, n13082, n13083, n13084, n13085,
         n13086, n13087, n13088, n13089, n13090, n13091, n13092, n13093,
         n13094, n13095, n13096, n13097, n13098, n13099, n13100, n13101,
         n13102, n13103, n13104, n13105, n13106, n13107, n13108, n13109,
         n13110, n13111, n13112, n13113, n13114, n13115, n13116, n13117,
         n13118, n13119, n13120, n13121, n13122, n13123, n13124, n13125,
         n13126, n13127, n13128, n13129, n13130, n13131, n13132, n13133,
         n13134, n13135, n13136, n13137, n13138, n13139, n13140, n13141,
         n13142, n13143, n13144, n13145, n13146, n13147, n13148, n13149,
         n13150, n13151, n13152, n13153, n13154, n13155, n13156, n13157,
         n13158, n13159, n13160, n13161, n13162, n13163, n13164, n13165,
         n13166, n13167, n13168, n13169, n13170, n13171, n13172, n13173,
         n13174, n13175, n13176, n13177, n13178, n13179, n13180, n13181,
         n13182, n13183, n13184, n13185, n13186, n13187, n13188, n13189,
         n13190, n13191, n13192, n13193, n13194, n13195, n13196, n13197,
         n13198, n13199, n13200, n13201, n13202, n13203, n13204, n13205,
         n13206, n13207, n13208, n13209, n13210, n13211, n13212, n13213,
         n13214, n13215, n13216, n13217, n13218, n13219, n13220, n13221,
         n13222, n13223, n13224, n13225, n13226, n13227, n13228, n13229,
         n13230, n13231, n13232, n13233, n13234, n13235, n13236, n13237,
         n13238, n13239, n13240, n13241, n13242, n13243, n13244, n13245,
         n13246, n13247, n13248, n13249, n13250, n13251, n13252, n13253,
         n13254, n13255, n13256, n13257, n13258, n13259, n13260, n13261,
         n13262, n13263, n13264, n13265, n13266, n13267, n13268, n13269,
         n13270, n13271, n13272, n13273, n13274, n13275, n13276, n13277,
         n13278, n13279, n13280, n13281, n13282, n13283, n13284, n13285,
         n13286, n13287, n13288, n13289, n13290, n13291, n13292, n13293,
         n13294, n13295, n13296, n13297, n13298, n13299, n13300, n13301,
         n13302, n13303, n13304, n13305, n13306, n13307, n13308, n13309,
         n13310, n13311, n13312, n13313, n13314, n13315, n13316, n13317,
         n13318, n13319, n13320, n13321, n13322, n13323, n13324, n13325,
         n13326, n13327, n13328, n13329, n13330, n13331, n13332, n13333,
         n13334, n13335, n13336, n13337, n13338, n13339, n13340, n13341,
         n13342, n13343, n13344, n13345, n13346, n13347, n13348, n13349,
         n13350, n13351, n13352, n13353, n13354, n13355, n13356, n13357,
         n13358, n13359, n13360, n13361, n13362, n13363, n13364, n13365,
         n13366, n13367, n13368, n13369, n13370, n13371, n13372, n13373,
         n13374, n13375, n13376, n13377, n13378, n13379, n13380, n13381,
         n13382, n13383, n13384, n13385, n13386, n13387, n13388, n13389,
         n13390, n13391, n13392, n13393, n13394, n13395, n13396, n13397,
         n13398, n13399, n13400, n13401, n13402, n13403, n13404, n13405,
         n13406, n13407, n13408, n13409, n13410, n13411, n13412, n13413,
         n13414, n13415, n13416, n13417, n13418, n13419, n13420, n13421,
         n13422, n13423, n13424, n13425, n13426, n13427, n13428, n13429,
         n13430, n13431, n13432, n13433, n13434, n13435, n13436, n13437,
         n13438, n13439, n13440, n13441, n13442, n13443, n13444, n13445,
         n13446, n13447, n13448, n13449, n13450, n13451, n13452, n13453,
         n13454, n13455, n13456, n13457, n13458, n13459, n13460, n13461,
         n13462, n13463, n13464, n13465, n13466, n13467, n13468, n13469,
         n13470, n13471, n13472, n13473, n13474, n13475, n13476, n13477,
         n13478, n13479, n13480, n13481, n13482, n13483, n13484, n13485,
         n13486, n13487, n13488, n13489, n13490, n13491, n13492, n13493,
         n13494, n13495, n13496, n13497, n13498, n13499, n13500, n13501,
         n13502, n13503, n13504, n13505, n13506, n13507, n13508, n13509,
         n13510, n13511, n13512, n13513, n13514, n13515, n13516, n13517,
         n13518, n13519, n13520, n13521, n13522, n13523, n13524, n13525,
         n13526, n13527, n13528, n13529, n13530, n13531, n13532, n13533,
         n13534, n13535, n13536, n13537, n13538, n13539, n13540, n13541,
         n13542, n13543, n13544, n13545, n13546, n13547, n13548, n13549,
         n13550, n13551, n13552, n13553, n13554, n13555, n13556, n13557,
         n13558, n13559, n13560, n13561, n13562, n13563, n13564, n13565,
         n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573,
         n13574, n13575, n13576, n13577, n13578, n13579, n13580, n13581,
         n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13589,
         n13590, n13591, n13592, n13593, n13594, n13595, n13596, n13597,
         n13598, n13599, n13600, n13601, n13602, n13603, n13604, n13605,
         n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613,
         n13614, n13615, n13616, n13617, n13618, n13619, n13620, n13621,
         n13622, n13623, n13624, n13625, n13626, n13627, n13628, n13629,
         n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13639,
         n13640, n13641, n13642, n13643, n13645, n13646, n13647, n13648,
         n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656,
         n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664,
         n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672,
         n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,
         n13682, n13683, n13684, n13686, n13687, n13688, n13689, intadd_8_A_5_,
         intadd_8_A_4_, intadd_8_A_3_, intadd_8_A_2_, intadd_8_B_6_,
         intadd_8_B_5_, intadd_8_B_4_, intadd_8_B_3_, intadd_8_B_2_,
         intadd_8_B_1_, intadd_8_n7, intadd_8_n6, intadd_8_n5, intadd_8_n4,
         intadd_8_n3, intadd_8_n2, intadd_8_n1, mult_x_433_n51, mult_x_433_n42,
         mult_x_433_n33, mult_x_433_n28, mult_x_433_n14, mult_x_433_n13,
         mult_x_433_n12, mult_x_433_n11, mult_x_433_n10, mult_x_433_n9,
         mult_x_433_n8, mult_x_433_n7, mult_x_433_n6, mult_x_433_n5,
         mult_x_431_n48, mult_x_431_n39, mult_x_431_n11, mult_x_431_n10,
         mult_x_431_n9, mult_x_431_n8, mult_x_431_n7, n13765, n13766, n13767,
         n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775,
         n13776, n13777, n13778, n13779, n13780, n13781, n13782, n13783,
         n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791,
         n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799,
         n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807,
         n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815,
         n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823,
         n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831,
         n13832, n13833, n13834, n13835, n13836, n13837, n13838, n13839,
         n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847,
         n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855,
         n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863,
         n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871,
         n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879,
         n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887,
         n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895,
         n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903,
         n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911,
         n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919,
         n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927,
         n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935,
         n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943,
         n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951,
         n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959,
         n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967,
         n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975,
         n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983,
         n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991,
         n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999,
         n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007,
         n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015,
         n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023,
         n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031,
         n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039,
         n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047,
         n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055,
         n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063,
         n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071,
         n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14079,
         n14080, n14081, n14082, n14083, n14084, n14085, n14086, n14087,
         n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095,
         n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103,
         n14104, n14105, n14106, n14107, n14108, n14109, n14110, n14111,
         n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119,
         n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127,
         n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135,
         n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143,
         n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151,
         n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14159,
         n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167,
         n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175,
         n14176, n14177, n14178, n14179, n14180, n14181, n14182, n14183,
         n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191,
         n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199,
         n14200, n14201, n14202, n14203, n14204, n14205, n14206, n14207,
         n14208, n14209, n14210, n14211, n14212, n14213, n14214, n14215,
         n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223,
         n14224, n14225, n14226, n14227, n14228, n14229, n14230, n14231,
         n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239,
         n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247,
         n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255,
         n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263,
         n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271,
         n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279,
         n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287,
         n14288, n14289, n14290, n14291, n14292, n14293, n14294, n14295,
         n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14303,
         n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311,
         n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319,
         n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327,
         n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335,
         n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343,
         n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351,
         n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359,
         n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367,
         n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375,
         n14376, n14377, n14378, n14379, n14380, n14381, n14382, n14383,
         n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391,
         n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399,
         n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407,
         n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415,
         n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423,
         n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431,
         n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439,
         n14440, n14441, n14442, n14443, n14444, n14445, n14446, n14447,
         n14448, n14449, n14450, n14451, n14452, n14453, n14454, n14455,
         n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14463,
         n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471,
         n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479,
         n14480, n14481, n14482, n14483, n14484, n14485, n14486, n14487,
         n14488, n14489, n14490, n14491, n14492, n14493, n14494, n14495,
         n14496, n14497, n14498, n14499, n14500, n14501, n14502, n14503,
         n14504, n14505, n14506, n14507, n14508, n14509, n14510, n14511,
         n14512, n14513, n14514, n14515, n14516, n14517, n14518, n14519,
         n14520, n14521, n14522, n14523, n14524, n14525, n14526, n14527,
         n14528, n14529, n14530, n14531, n14532, n14533, n14534, n14535,
         n14536, n14537, n14538, n14539, n14540, n14541, n14542, n14543,
         n14544, n14545, n14546, n14547, n14548, n14549, n14550, n14551,
         n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559,
         n14560, n14561, n14562, n14563, n14564, n14565, n14566, n14567,
         n14568, n14569, n14570, n14571, n14572, n14573, n14574, n14575,
         n14576, n14577, n14578, n14579, n14580, n14581, n14582, n14583,
         n14584, n14585, n14586, n14587, n14588, n14589, n14590, n14591,
         n14592, n14593, n14594, n14595, n14596, n14597, n14598, n14599,
         n14600, n14601, n14602, n14603, n14604, n14605, n14606, n14607,
         n14608, n14609, n14610, n14611, n14612, n14613, n14614, n14615,
         n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623,
         n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631,
         n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639,
         n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647,
         n14648, n14649, n14650, n14651, n14652, n14653, n14654, n14655,
         n14656, n14657, n14658, n14659, n14660, n14661, n14662, n14663,
         n14664, n14665, n14666, n14667, n14668, n14669, n14670, n14671,
         n14672, n14673, n14674, n14675, n14676, n14677, n14678, n14679,
         n14680, n14681, n14682, n14683, n14684, n14685, n14686, n14687,
         n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695,
         n14696, n14697, n14698, n14699, n14700, n14701, n14702, n14703,
         n14704, n14705, n14706, n14707, n14708, n14709, n14710, n14711,
         n14712, n14713, n14714, n14715, n14716, n14717, n14718, n14719,
         n14720, n14721, n14722, n14723, n14724, n14725, n14726, n14727,
         n14728, n14729, n14730, n14731, n14732, n14733, n14734, n14735,
         n14736, n14737, n14738, n14739, n14740, n14741, n14742, n14743,
         n14744, n14745, n14746, n14747, n14748, n14749, n14750, n14751,
         n14752, n14753, n14754, n14755, n14756, n14757, n14758, n14759,
         n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14767,
         n14768, n14769, n14770, n14771, n14772, n14773, n14774, n14775,
         n14776, n14777, n14778, n14779, n14780, n14781, n14782, n14783,
         n14784, n14785, n14786, n14787, n14788, n14789, n14790, n14791,
         n14792, n14793, n14794, n14795, n14796, n14797, n14798, n14799,
         n14800, n14801, n14802, n14803, n14804, n14805, n14806, n14807,
         n14808, n14809, n14810, n14811, n14812, n14813, n14814, n14815,
         n14816, n14817, n14818, n14819, n14820, n14821, n14822, n14823,
         n14824, n14825, n14826, n14827, n14828, n14829, n14830, n14831,
         n14832, n14833, n14834, n14835, n14836, n14837, n14838, n14839,
         n14840, n14841, n14842, n14843, n14844, n14845, n14846, n14847,
         n14848, n14849, n14850, n14851, n14852, n14853, n14854, n14855,
         n14856, n14857, n14858, n14859, n14860, n14861, n14862, n14863,
         n14864, n14865, n14866, n14867, n14868, n14869, n14870, n14871,
         n14872, n14873, n14874, n14875, n14876, n14877, n14878, n14879,
         n14880, n14881, n14882, n14883, n14884, n14885, n14886, n14887,
         n14888, n14889, n14890, n14891, n14892, n14893, n14894, n14895,
         n14896, n14897, n14898, n14899, n14900, n14901, n14902, n14903,
         n14904, n14905, n14906, n14907, n14908, n14909, n14910, n14911,
         n14912, n14913, n14914, n14915, n14916, n14917, n14918, n14919,
         n14920, n14921, n14922, n14923, n14924, n14925, n14926, n14927,
         n14928, n14929, n14930, n14931, n14932, n14933, n14934, n14935,
         n14936, n14937, n14938, n14939, n14940, n14941, n14942, n14943,
         n14944, n14945, n14946, n14947, n14948, n14949, n14950, n14951,
         n14952, n14953, n14954, n14955, n14956, n14957, n14958, n14959,
         n14960, n14961, n14962, n14963, n14964, n14965, n14966, n14967,
         n14968, n14969, n14970, n14971, n14972, n14973, n14974, n14975,
         n14976, n14977, n14978, n14979, n14980, n14981, n14982, n14983,
         n14984, n14985, n14986, n14987, n14988, n14989, n14990, n14991,
         n14992, n14993, n14994, n14995, n14996, n14997, n14998, n14999,
         n15000, n15001, n15002, n15003, n15004, n15005, n15006, n15007,
         n15008, n15009, n15010, n15011, n15012, n15013, n15014, n15015,
         n15016, n15017, n15018, n15019, n15020, n15021, n15022, n15023,
         n15024, n15025, n15026, n15027, n15028, n15029, n15030, n15031,
         n15032, n15033, n15034, n15035, n15036, n15037, n15038, n15039,
         n15040, n15041, n15042, n15043, n15044, n15045, n15046, n15047,
         n15048, n15049, n15050, n15051, n15052, n15053, n15054, n15055,
         n15056, n15057, n15058, n15059, n15060, n15061, n15062, n15063,
         n15064, n15065, n15066, n15067, n15068, n15069, n15070, n15071,
         n15072, n15073, n15074, n15075, n15076, n15077, n15078, n15079,
         n15080, n15081, n15082, n15083, n15084, n15085, n15086, n15087,
         n15088, n15089, n15090, n15091, n15092, n15093, n15094, n15095,
         n15096, n15097, n15098, n15099, n15100, n15101, n15102, n15103,
         n15104, n15105, n15106, n15107, n15108, n15109, n15110, n15111,
         n15112, n15113, n15114, n15115, n15116, n15117, n15118, n15119,
         n15120, n15121, n15122, n15123, n15124, n15125, n15126, n15127,
         n15128, n15129, n15130, n15131, n15132, n15133, n15134, n15135,
         n15136, n15137, n15138, n15139, n15140, n15141, n15142, n15143,
         n15144, n15145, n15146, n15147, n15148, n15149, n15150, n15151,
         n15152, n15153, n15154, n15155, n15156, n15157, n15158, n15159,
         n15160, n15161, n15162, n15163, n15164, n15165, n15166, n15167,
         n15168, n15169, n15170, n15171, n15172, n15173, n15174, n15175,
         n15176, n15177, n15178, n15179, n15180, n15181, n15182, n15183,
         n15184, n15185, n15186, n15187, n15188, n15189, n15190, n15191,
         n15192, n15193, n15194, n15195, n15196, n15197, n15198, n15199,
         n15200, n15201, n15202, n15203, n15204, n15205, n15206, n15207,
         n15208, n15209, n15210, n15211, n15212, n15213, n15214, n15215,
         n15216, n15217, n15218, n15219, n15220, n15221, n15222, n15223,
         n15224, n15225, n15226, n15227, n15228, n15229, n15230, n15231,
         n15232, n15233, n15234, n15235, n15236, n15237, n15238, n15239,
         n15240, n15241, n15242, n15243, n15244, n15245, n15246, n15247,
         n15248, n15249, n15250, n15251, n15252, n15253, n15254, n15255,
         n15256, n15257, n15258, n15259, n15260, n15261, n15262, n15263,
         n15264, n15265, n15266, n15267, n15268, n15269, n15270, n15271,
         n15272, n15273, n15274, n15275, n15276, n15277, n15278, n15279,
         n15280, n15281, n15282, n15283, n15284, n15285, n15286, n15287,
         n15288, n15289, n15290, n15291, n15292, n15293, n15294, n15295,
         n15296, n15297, n15298, n15299, n15300, n15301, n15302, n15303,
         n15304, n15305, n15306, n15307, n15308, n15309, n15310, n15311,
         n15312, n15313, n15314, n15315, n15316, n15317, n15318, n15319,
         n15320, n15321, n15322, n15323, n15324, n15325, n15326, n15327,
         n15328, n15329, n15330, n15331, n15332, n15333, n15334, n15335,
         n15336, n15337, n15338, n15339, n15340, n15341, n15342, n15343,
         n15344, n15345, n15346, n15347, n15348, n15349, n15350, n15351,
         n15352, n15353, n15354, n15355, n15356, n15357, n15358, n15359,
         n15360, n15361, n15362, n15363, n15364, n15365, n15366, n15367,
         n15368, n15369, n15370, n15371, n15372, n15373, n15374, n15375,
         n15376, n15377, n15378, n15379, n15380, n15381, n15382, n15383,
         n15384, n15385, n15386, n15387, n15388, n15389, n15390, n15391,
         n15392, n15393, n15394, n15395, n15396, n15397, n15398, n15399,
         n15400, n15401, n15402, n15403, n15404, n15405, n15406, n15407,
         n15408, n15409, n15410, n15411, n15412, n15413, n15414, n15415,
         n15416, n15417, n15418, n15419, n15420, n15421, n15422, n15423,
         n15424, n15425, n15426, n15427, n15428, n15429, n15430, n15431,
         n15432, n15433, n15434, n15435, n15436, n15437, n15438, n15439,
         n15440, n15441, n15442, n15443, n15444, n15445, n15446, n15447,
         n15448, n15449, n15450, n15451, n15452, n15453, n15454, n15455,
         n15456, n15457, n15458, n15459, n15460, n15461, n15462, n15463,
         n15464, n15465, n15466, n15467, n15468, n15469, n15470, n15471,
         n15472, n15473, n15474, n15475, n15476, n15477, n15478, n15479,
         n15480, n15481, n15482, n15483, n15484, n15485, n15486, n15487,
         n15488, n15489, n15490, n15491, n15492, n15493, n15494, n15495,
         n15496, n15497, n15498, n15499, n15500, n15501, n15502, n15503,
         n15504, n15505, n15506, n15507, n15508, n15509, n15510, n15511,
         n15512, n15513, n15514, n15515, n15516, n15517, n15518, n15519,
         n15520, n15521, n15522, n15523, n15524, n15525, n15526, n15527,
         n15528, n15529, n15530, n15531, n15532, n15533, n15534, n15535,
         n15536, n15537, n15538, n15539, n15540, n15541, n15542, n15543,
         n15544, n15545, n15546, n15547, n15548, n15549, n15550, n15551,
         n15552, n15553, n15554, n15555, n15556, n15557, n15558, n15559,
         n15560, n15561, n15562, n15563, n15564, n15565, n15566, n15567,
         n15568, n15569, n15570, n15571, n15572, n15573, n15574, n15575,
         n15576, n15577, n15578, n15579, n15580, n15581, n15582, n15583,
         n15584, n15585, n15586, n15587, n15588, n15589, n15590, n15591,
         n15592, n15593, n15594, n15595, n15596, n15597, n15598, n15599,
         n15600, n15601, n15602, n15603, n15604, n15605, n15606, n15607,
         n15608, n15609, n15610, n15611, n15612, n15613, n15614, n15615,
         n15616, n15617, n15618, n15619, n15620, n15621, n15622, n15623,
         n15624, n15625, n15626, n15627, n15628, n15629, n15630, n15631,
         n15632, n15633, n15634, n15635, n15636, n15637, n15638, n15639,
         n15640, n15641, n15642, n15643, n15644, n15645, n15646, n15647,
         n15648, n15649, n15650, n15651, n15652, n15653, n15654, n15655,
         n15656, n15657, n15658, n15659, n15660, n15661, n15662, n15663,
         n15664, n15665, n15666, n15667, n15668, n15669, n15670, n15671,
         n15672, n15673, n15674, n15675, n15676, n15677, n15678, n15679,
         n15680, n15681, n15682, n15683, n15684, n15685, n15686, n15687,
         n15688, n15689, n15690, n15691, n15692, n15693, n15694, n15695,
         n15696, n15697, n15698, n15699, n15700, n15701, n15702, n15703,
         n15704, n15705, n15706, n15707, n15708, n15709, n15710, n15711,
         n15712, n15713, n15714, n15715, n15716, n15717, n15718, n15719,
         n15720, n15721, n15722, n15723, n15724, n15725, n15726, n15727,
         n15728, n15729, n15730, n15731, n15732, n15733, n15734, n15735,
         n15736, n15737, n15738, n15739, n15740, n15741, n15742, n15743,
         n15744, n15745, n15746, n15747, n15748, n15749, n15750, n15751,
         n15752, n15753, n15754, n15755, n15756, n15757, n15758, n15759,
         n15760, n15761, n15762, n15763, n15764, n15765, n15766, n15767,
         n15768, n15769, n15770, n15771, n15772, n15773, n15774, n15775,
         n15776, n15777, n15778, n15779, n15780, n15781, n15782, n15783,
         n15784, n15785, n15786, n15787, n15788, n15789, n15790, n15791,
         n15792, n15793, n15794, n15795, n15796, n15797, n15798, n15799,
         n15800, n15801, n15802, n15803, n15804, n15805, n15806, n15807,
         n15808, n15809, n15810, n15811, n15812, n15813, n15814, n15815,
         n15816, n15817, n15818, n15819, n15820, n15821, n15822, n15823,
         n15824, n15825, n15826, n15827, n15828, n15829, n15830, n15831,
         n15832, n15833, n15834, n15835, n15836, n15837, n15838, n15839,
         n15840, n15841, n15842, n15843, n15844, n15845, n15846, n15847,
         n15848, n15849, n15850, n15851, n15852, n15853, n15854, n15855,
         n15856, n15857, n15858, n15859, n15860, n15861, n15862, n15863,
         n15864, n15865, n15866, n15867, n15868, n15869, n15870, n15871,
         n15872, n15873, n15874, n15875, n15876, n15877, n15878, n15879,
         n15880, n15881, n15882, n15883, n15884, n15885, n15886, n15887,
         n15888, n15889, n15890, n15891, n15892, n15893, n15894, n15895,
         n15896, n15897, n15898, n15899, n15900, n15901, n15902, n15903,
         n15904, n15905, n15906, n15907, n15908, n15909, n15910, n15911,
         n15912, n15913, n15914, n15915, n15916, n15917, n15918, n15919,
         n15920, n15921, n15922, n15923, n15924, n15925, n15926, n15927,
         n15928, n15929, n15930, n15931, n15932, n15933, n15934, n15935,
         n15936, n15937, n15938, n15939, n15940, n15941, n15942, n15943,
         n15944, n15945, n15946, n15947, n15948, n15949, n15950, n15951,
         n15952, n15953, n15954, n15955, n15956, n15957, n15958, n15959,
         n15960, n15961, n15962, n15963, n15964, n15965, n15966, n15967,
         n15968, n15969, n15970, n15971, n15972, n15973, n15974, n15975,
         n15976, n15977, n15978, n15979, n15980, n15981, n15982, n15983,
         n15984, n15985, n15986, n15987, n15988, n15989, n15990, n15991,
         n15992, n15993, n15994, n15995, n15996, n15997, n15998, n15999,
         n16000, n16001, n16002, n16003, n16004, n16005, n16006, n16007,
         n16008, n16009, n16010, n16011, n16012, n16013, n16014, n16015,
         n16016, n16017, n16018, n16019, n16020, n16021, n16022, n16023,
         n16024, n16025, n16026, n16027, n16028, n16029, n16030, n16031,
         n16032, n16033, n16034, n16035, n16036, n16037, n16038, n16039,
         n16040, n16041, n16042, n16043, n16044, n16045, n16046, n16047,
         n16048, n16049, n16050, n16051, n16052, n16053, n16054, n16055,
         n16056, n16057, n16058, n16059, n16060, n16061, n16062, n16063,
         n16064, n16065, n16066, n16067, n16068, n16069, n16070, n16071,
         n16072, n16073, n16074, n16075, n16076, n16077, n16078, n16079,
         n16080, n16081, n16082, n16083, n16084, n16085, n16086, n16087,
         n16088, n16089, n16090, n16091, n16092, n16093, n16094, n16095,
         n16096, n16097, n16098, n16099, n16100, n16101, n16102, n16103,
         n16104, n16105, n16106, n16107, n16108, n16109, n16110, n16111,
         n16112, n16113, n16114, n16115, n16116, n16117, n16118, n16119,
         n16120, n16121, n16122, n16123, n16124, n16125, n16126, n16127,
         n16128, n16129, n16130, n16131, n16132, n16133, n16134, n16135,
         n16136, n16137, n16138, n16139, n16140, n16141, n16142, n16143,
         n16144, n16145, n16146, n16147, n16148, n16149, n16150, n16151,
         n16152, n16153, n16154, n16155, n16156, n16157, n16158, n16159,
         n16160, n16161, n16162, n16163, n16164, n16165, n16166, n16167,
         n16168, n16169, n16170, n16171, n16172, n16173, n16174, n16175,
         n16176, n16177, n16178, n16179, n16180, n16181, n16182, n16183,
         n16184, n16185, n16186, n16187, n16188, n16189, n16190, n16191,
         n16192, n16193, n16194, n16195, n16196, n16197, n16198, n16199,
         n16200, n16201, n16202, n16203, n16204, n16205, n16206, n16207,
         n16208, n16209, n16210, n16211, n16212, n16213, n16214, n16215,
         n16216, n16217, n16218, n16219, n16220, n16221, n16222, n16223,
         n16224, n16225, n16226, n16227, n16228, n16229, n16230, n16231,
         n16232, n16233, n16234, n16235, n16236, n16237, n16238, n16239,
         n16240, n16241, n16242, n16243, n16244, n16245, n16246, n16247,
         n16248, n16249, n16250, n16251, n16252, n16253, n16254, n16255,
         n16256, n16257, n16258, n16259, n16260, n16261, n16262, n16263,
         n16264, n16265, n16266, n16267, n16268, n16269, n16270, n16271,
         n16272, n16273, n16274, n16275, n16276, n16277, n16278, n16279,
         n16280, n16281, n16282, n16283, n16284, n16285, n16286, n16287,
         n16288, n16289, n16290, n16291, n16292, n16293, n16294, n16295,
         n16296, n16297, n16298, n16299, n16300, n16301, n16302, n16303,
         n16304, n16305, n16306, n16307, n16308, n16309, n16310, n16311,
         n16312, n16313, n16314, n16315, n16316, n16317, n16318, n16319,
         n16320, n16321, n16322, n16323, n16324, n16325, n16326, n16327,
         n16328, n16329, n16330, n16331, n16332, n16333, n16334, n16335,
         n16336, n16337, n16338, n16339, n16340, n16341, n16342, n16343,
         n16344, n16345, n16346, n16347, n16348, n16349, n16350, n16351,
         n16352, n16353, n16354, n16355, n16356, n16357, n16358, n16359,
         n16360, n16361, n16362, n16363, n16364, n16365, n16366, n16367,
         n16368, n16369, n16370, n16371, n16372, n16373, n16374, n16375,
         n16376, n16377, n16378, n16379, n16380, n16381, n16382, n16383,
         n16384, n16385, n16386, n16387, n16388, n16389, n16390, n16391,
         n16392, n16393, n16394, n16395, n16396, n16397, n16398, n16399,
         n16400, n16401, n16402, n16403, n16404, n16405, n16406, n16407,
         n16408, n16409, n16410, n16411, n16412, n16413, n16414, n16415,
         n16416, n16417, n16418, n16419, n16420, n16421, n16422, n16423,
         n16424, n16425, n16426, n16427, n16428, n16429, n16430, n16431,
         n16432, n16433, n16434, n16435, n16436, n16437, n16438, n16439,
         n16440, n16441, n16442, n16443, n16444, n16445, n16446, n16447,
         n16448, n16449, n16450, n16451, n16452, n16453, n16454, n16455,
         n16456, n16457, n16458, n16459, n16460, n16461, n16462, n16463,
         n16464, n16465, n16466, n16467, n16468, n16469, n16470, n16471,
         n16472, n16473, n16474, n16475, n16476, n16477, n16478, n16479,
         n16480, n16481, n16482, n16483, n16484, n16485, n16486, n16487,
         n16488, n16489, n16490, n16491, n16492, n16493, n16494, n16495,
         n16496, n16497, n16498, n16499, n16500, n16501, n16502, n16503,
         n16504, n16505, n16506, n16507, n16508, n16509, n16510, n16511,
         n16512, n16513, n16514, n16515, n16516, n16517, n16518, n16519,
         n16520, n16521, n16522, n16523, n16524, n16525, n16526, n16527,
         n16528, n16529, n16530, n16531, n16532, n16533, n16534, n16535,
         n16536, n16537, n16538, n16539, n16540, n16541, n16542, n16543,
         n16544, n16545, n16546, n16547, n16548, n16549, n16550, n16551,
         n16552, n16553, n16554, n16555, n16556, n16557, n16558, n16559,
         n16560, n16561, n16562, n16563, n16564, n16565, n16566, n16567,
         n16568, n16569, n16570, n16571, n16572, n16573, n16574, n16575,
         n16576, n16577, n16578, n16579, n16580, n16581, n16582, n16583,
         n16584, n16585, n16586, n16587, n16588, n16589, n16590, n16591,
         n16592, n16593, n16594, n16595, n16596, n16597, n16598, n16599,
         n16600, n16601, n16602, n16603, n16604, n16605, n16606, n16607,
         n16608, n16609, n16610, n16611, n16612, n16613, n16614, n16615,
         n16616, n16617, n16618, n16619, n16620, n16621, n16622, n16623,
         n16624, n16625, n16626, n16627, n16628, n16629, n16630, n16631,
         n16632, n16633, n16634, n16635, n16636, n16637, n16638, n16639,
         n16640, n16641, n16642, n16643, n16644, n16645, n16646, n16647,
         n16648, n16649, n16650, n16651, n16652, n16653, n16654, n16655,
         n16656, n16657, n16658, n16659, n16660, n16661, n16662, n16663,
         n16664, n16665, n16666, n16667, n16668, n16669, n16670, n16671,
         n16672, n16673, n16674, n16675, n16676, n16677, n16678, n16679,
         n16680, n16681, n16682, n16683, n16684, n16685, n16686, n16687,
         n16688, n16689, n16690, n16691, n16692, n16693, n16694, n16695,
         n16696, n16697, n16698, n16699, n16700, n16701, n16702, n16703,
         n16704, n16705, n16706, n16707, n16708, n16709, n16710, n16711,
         n16712, n16713, n16714, n16715, n16716, n16717, n16718, n16719,
         n16720, n16721, n16722, n16723, n16724, n16725, n16726, n16727,
         n16728, n16729, n16730, n16731, n16732, n16733, n16734, n16735,
         n16736, n16737, n16738, n16739, n16740, n16741, n16742, n16743,
         n16744, n16745, n16746, n16747, n16748, n16749, n16750, n16751,
         n16752, n16753, n16754, n16755, n16756, n16757, n16758, n16759,
         n16760, n16761, n16762, n16763, n16764, n16765, n16766, n16767,
         n16768, n16769, n16770, n16771, n16772, n16773, n16774, n16775,
         n16776, n16777, n16778, n16779, n16780, n16781, n16782, n16783,
         n16784, n16785, n16786, n16787, n16788, n16789, n16790, n16791,
         n16792, n16793, n16794, n16795, n16796, n16797, n16798, n16799,
         n16800, n16801, n16802, n16803, n16804, n16805, n16806, n16807,
         n16808, n16809, n16810, n16811, n16812, n16813, n16814, n16815,
         n16816, n16817, n16818, n16819, n16820, n16821, n16822, n16823,
         n16824, n16825, n16826, n16827, n16828, n16829, n16830, n16831,
         n16832, n16833, n16834, n16835, n16836, n16837, n16838, n16839,
         n16840, n16841, n16842, n16843, n16844, n16845, n16846, n16847,
         n16848, n16849, n16850, n16851, n16852, n16853, n16854, n16855,
         n16856, n16857, n16858, n16859, n16860, n16861, n16862, n16863,
         n16864, n16865, n16866, n16867, n16868, n16869, n16870, n16871,
         n16872, n16873, n16874, n16875, n16876, n16877, n16878, n16879,
         n16880, n16881, n16882, n16883, n16884, n16885, n16886, n16887,
         n16888, n16889, n16890, n16891, n16892, n16893, n16894, n16895,
         n16896, n16897, n16898, n16899, n16900, n16901, n16902, n16903,
         n16904, n16905, n16906, n16907, n16908, n16909, n16910, n16911,
         n16912, n16913, n16914, n16915, n16916, n16917, n16918, n16919,
         n16920, n16921, n16922, n16923, n16924, n16925, n16926, n16927,
         n16928, n16929, n16930, n16931, n16932, n16933, n16934, n16935,
         n16936, n16937, n16938, n16939, n16940, n16941, n16942, n16943,
         n16944, n16945, n16946, n16947, n16948, n16949, n16950, n16951,
         n16952, n16953, n16954, n16955, n16956, n16957, n16958, n16959,
         n16960, n16961, n16962, n16963, n16964, n16965, n16966, n16967,
         n16968, n16969, n16970, n16971, n16972, n16973, n16974, n16975,
         n16976, n16977, n16978, n16979, n16980, n16981, n16982, n16983,
         n16984, n16985, n16986, n16987, n16988, n16989, n16990, n16991,
         n16992, n16993, n16994, n16995, n16996, n16997, n16998, n16999,
         n17000, n17001, n17002, n17003, n17004, n17005, n17006, n17007,
         n17008, n17009, n17010, n17011, n17012, n17013, n17014, n17015,
         n17016, n17017, n17018, n17019, n17020, n17021, n17022, n17023,
         n17024, n17025, n17026, n17027, n17028, n17029, n17030, n17031,
         n17032, n17033, n17034, n17035, n17036, n17037, n17038, n17039,
         n17040, n17041, n17042, n17043, n17044, n17045, n17046, n17047,
         n17048, n17049, n17050, n17051, n17052, n17053, n17054, n17055,
         n17056, n17057, n17058, n17059, n17060, n17061, n17062, n17063,
         n17064, n17065, n17066, n17067, n17068, n17069, n17070, n17071,
         n17072, n17073, n17074, n17075, n17076, n17077, n17078, n17079,
         n17080, n17081, n17082, n17083, n17084, n17085, n17086, n17087,
         n17088, n17089, n17090, n17091, n17092, n17093, n17094, n17095,
         n17096, n17097, n17098, n17099, n17100, n17101, n17102, n17103,
         n17104, n17105, n17106, n17107, n17108, n17109, n17110, n17111,
         n17112, n17113, n17114, n17115, n17116, n17117, n17118, n17119,
         n17120, n17121, n17122, n17123, n17124, n17125, n17126, n17127,
         n17128, n17129, n17130, n17131, n17132, n17133, n17134, n17135,
         n17136, n17137, n17138, n17139, n17140, n17141, n17142, n17143,
         n17144, n17145, n17146, n17147, n17148, n17149, n17150, n17151,
         n17152, n17153, n17154, n17155, n17156, n17157, n17158, n17159,
         n17160, n17161, n17162, n17163, n17164, n17165, n17166, n17167,
         n17168, n17169, n17170, n17171, n17172, n17173, n17174, n17175,
         n17176, n17177, n17178, n17179, n17180, n17181, n17182, n17183,
         n17184, n17185, n17186, n17187, n17188, n17189, n17190, n17191,
         n17192, n17193, n17194, n17195, n17196, n17197, n17198, n17199,
         n17200, n17201, n17202, n17203, n17204, n17205, n17206, n17207,
         n17208, n17209, n17210, n17211, n17212, n17213, n17214, n17215,
         n17216, n17217, n17218, n17219, n17220, n17221, n17222, n17223,
         n17224, n17225, n17226, n17227, n17228, n17229, n17230, n17231,
         n17232, n17233, n17234, n17235, n17236, n17237, n17238, n17239,
         n17240, n17241, n17242, n17243, n17244, n17245, n17246, n17247,
         n17248, n17249, n17250, n17251, n17252, n17253, n17254, n17255,
         n17256, n17257, n17258, n17259, n17260, n17261, n17262, n17263,
         n17264, n17265, n17266, n17267, n17268, n17269, n17270, n17271,
         n17272, n17273, n17274, n17275, n17276, n17277, n17278, n17279,
         n17280, n17281, n17282, n17283, n17284, n17285, n17286, n17287,
         n17288, n17289, n17290, n17291, n17292, n17293, n17294, n17295,
         n17296, n17297, n17298, n17299, n17300, n17301, n17302, n17303,
         n17304, n17305, n17306, n17307, n17308, n17309, n17310, n17311,
         n17312, n17313, n17314, n17315, n17316, n17317, n17318, n17319,
         n17320, n17321, n17322, n17323, n17324, n17325, n17326, n17327,
         n17328, n17329, n17330, n17331, n17332, n17333, n17334, n17335,
         n17336, n17337, n17338, n17339, n17340, n17341, n17342, n17343,
         n17344, n17345, n17346, n17347, n17348, n17349, n17350, n17351,
         n17352, n17353, n17354, n17355, n17356, n17357, n17358, n17359,
         n17360, n17361, n17362, n17363, n17364, n17365, n17366, n17367,
         n17368, n17369, n17370, n17371, n17372, n17373, n17374, n17375,
         n17376, n17377, n17378, n17379, n17380, n17381, n17382, n17383,
         n17384, n17385, n17386, n17387, n17388, n17389, n17390, n17391,
         n17392, n17393, n17394, n17395, n17396, n17397, n17398, n17399,
         n17400, n17401, n17402, n17403, n17404, n17405, n17406, n17407,
         n17408, n17409, n17410, n17411, n17412, n17413, n17414, n17415,
         n17416, n17417, n17418, n17419, n17420, n17421, n17422, n17423,
         n17424, n17425, n17426, n17427, n17428, n17429, n17430, n17431,
         n17432, n17433, n17434, n17435, n17436, n17437, n17438, n17439,
         n17440, n17441, n17442, n17443, n17444, n17445, n17446, n17447,
         n17448, n17449, n17450, n17451, n17452, n17453, n17454, n17455,
         n17456, n17457, n17458, n17459, n17460, n17461, n17462, n17463,
         n17464, n17465, n17466, n17467, n17468, n17469, n17470, n17471,
         n17472, n17473, n17474, n17475, n17476, n17477, n17478, n17479,
         n17480, n17481, n17482, n17483, n17484, n17485, n17486, n17487,
         n17488, n17489, n17490, n17491, n17492, n17493, n17494, n17495,
         n17496, n17497, n17498, n17499, n17500, n17501, n17502, n17503,
         n17504, n17505, n17506, n17507, n17508, n17509, n17510, n17511,
         n17512, n17513, n17514, n17515, n17516, n17517, n17518, n17519,
         n17520, n17521, n17522, n17523, n17524, n17525, n17526, n17527,
         n17528, n17529, n17530, n17531, n17532, n17533, n17534, n17535,
         n17536, n17537, n17538, n17539, n17540, n17541, n17542, n17543,
         n17544, n17545, n17546, n17547, n17548, n17549, n17550, n17551,
         n17552, n17553, n17554, n17555, n17556, n17557, n17558, n17559,
         n17560, n17561, n17562, n17563, n17564, n17565, n17566, n17567,
         n17568, n17569, n17570, n17571, n17572, n17573, n17574, n17575,
         n17576, n17577, n17578, n17579, n17580, n17581, n17582, n17583,
         n17584, n17585, n17586, n17587, n17588, n17589, n17590, n17591,
         n17592, n17593, n17594, n17595, n17596, n17597, n17598, n17599,
         n17600, n17601, n17602, n17603, n17604, n17605, n17606, n17607,
         n17608, n17609, n17610, n17611, n17612, n17613, n17614, n17615,
         n17616, n17617, n17618, n17619, n17620, n17621, n17622, n17623,
         n17624, n17625, n17626, n17627, n17628, n17629, n17630, n17631,
         n17632, n17633, n17634, n17635, n17636, n17637, n17638, n17639,
         n17640, n17641, n17642, n17643, n17644, n17645, n17646, n17647,
         n17648, n17649, n17650, n17651, n17652, n17653, n17654, n17655,
         n17656, n17657, n17658, n17659, n17660, n17661, n17662, n17663,
         n17664, n17665, n17666, n17667, n17668, n17669, n17670, n17671,
         n17672, n17673, n17674, n17675, n17676, n17677, n17678, n17679,
         n17680, n17681, n17682, n17683, n17684, n17685, n17686, n17687,
         n17688, n17689, n17690, n17691, n17692, n17693, n17694, n17695,
         n17696, n17697, n17698, n17699, n17700, n17701, n17702, n17703,
         n17704, n17705, n17706, n17707, n17708, n17709, n17710, n17711,
         n17712, n17713, n17714, n17715, n17716, n17717, n17718, n17719,
         n17720, n17721, n17722, n17723, n17724, n17725, n17726, n17727,
         n17728, n17729, n17730, n17731, n17732, n17733, n17734, n17735,
         n17736, n17737, n17738, n17739, n17740, n17741, n17742, n17743,
         n17744, n17745, n17746, n17747, n17748, n17749, n17750, n17751,
         n17752, n17753, n17754, n17755, n17756, n17757, n17758, n17759,
         n17760, n17761, n17762, n17763, n17764, n17765, n17766, n17767,
         n17768, n17769, n17770, n17771, n17772, n17773, n17774, n17775,
         n17776, n17777, n17778, n17779, n17780, n17781, n17782, n17783,
         n17784, n17785, n17786, n17787, n17788, n17789, n17790, n17791,
         n17792, n17793, n17794, n17795, n17796, n17797, n17798, n17799,
         n17800, n17801, n17802, n17803, n17804, n17805, n17806, n17807,
         n17808, n17809, n17810, n17811, n17812, n17813, n17814, n17815,
         n17816, n17817, n17818, n17819, n17820, n17821, n17822, n17823,
         n17824, n17825, n17826, n17827, n17828, n17829, n17830, n17831,
         n17832, n17833, n17834, n17835, n17836, n17837, n17838, n17839,
         n17840, n17841, n17842, n17843, n17844, n17845, n17846, n17847,
         n17848, n17849, n17850, n17851, n17852, n17853, n17854, n17855,
         n17856, n17857, n17858, n17859, n17860, n17861, n17862, n17863,
         n17864, n17865, n17866, n17867, n17868, n17869, n17870, n17871,
         n17872, n17873, n17874, n17875, n17876, n17877, n17878, n17879,
         n17880, n17881, n17882, n17883, n17884, n17885, n17886, n17887,
         n17888, n17889, n17890, n17891, n17892, n17893, n17894, n17895,
         n17896, n17897, n17898, n17899, n17900, n17901, n17902, n17903,
         n17904, n17905, n17906, n17907, n17908, n17909, n17910, n17911,
         n17912, n17913, n17914, n17915, n17916, n17917, n17918, n17919,
         n17920, n17921, n17922, n17923, n17924, n17925, n17926, n17927,
         n17928, n17929, n17930, n17931, n17932, n17933, n17934, n17935,
         n17936, n17937, n17938, n17939, n17940, n17941, n17942, n17943,
         n17944, n17945, n17946, n17947, n17948, n17949, n17950, n17951,
         n17952, n17953, n17954, n17955, n17956, n17957, n17958, n17959,
         n17960, n17961, n17962, n17963, n17964, n17965, n17966, n17967,
         n17968, n17969, n17970, n17971, n17972, n17973, n17974, n17975,
         n17976, n17977, n17978, n17979, n17980, n17981, n17982, n17983,
         n17984, n17985, n17986, n17987, n17988, n17989, n17990, n17991,
         n17992, n17993, n17994, n17995, n17996, n17997, n17998, n17999,
         n18000, n18001, n18002, n18003, n18004, n18005, n18006, n18007,
         n18008, n18009, n18010, n18011, n18012, n18013, n18014, n18015,
         n18016, n18017, n18018, n18019, n18020, n18021, n18022, n18023,
         n18024, n18025, n18026, n18027, n18028, n18029, n18030, n18031,
         n18032, n18033, n18034, n18035, n18036, n18037, n18038, n18039,
         n18040, n18041, n18042, n18043, n18044, n18045, n18046, n18047,
         n18048, n18049, n18050, n18051, n18052, n18053, n18054, n18055,
         n18056, n18057, n18058, n18059, n18060, n18061, n18062, n18063,
         n18064, n18065, n18066, n18067, n18068, n18069, n18070, n18071,
         n18072, n18073, n18074, n18075, n18076, n18077, n18078, n18079,
         n18080, n18081, n18082, n18083, n18084, n18085, n18086, n18087,
         n18088, n18089, n18090, n18091, n18092, n18093, n18094, n18095,
         n18096, n18097, n18098, n18099, n18100, n18101, n18102, n18103,
         n18104, n18105, n18106, n18107, n18108, n18109, n18110, n18111,
         n18112, n18113, n18114, n18115, n18116, n18117, n18118, n18119,
         n18120, n18121, n18122, n18123, n18124, n18125, n18126, n18127,
         n18128, n18129, n18130, n18131, n18132, n18133, n18134, n18135,
         n18136, n18137, n18138, n18139, n18140, n18141, n18142, n18143,
         n18144, n18145, n18146, n18147, n18148, n18149, n18150, n18151,
         n18152, n18153, n18154, n18155, n18156, n18157, n18158, n18159,
         n18160, n18161, n18162, n18163, n18164, n18165, n18166, n18167,
         n18168, n18169, n18170, n18171, n18172, n18173, n18174, n18175,
         n18176, n18177, n18178, n18179, n18180, n18181, n18182, n18183,
         n18184, n18185, n18186, n18187, n18188, n18189, n18190, n18191,
         n18192, n18193, n18194, n18195, n18196, n18197, n18198, n18199,
         n18200, n18201, n18202, n18203, n18204, n18205, n18206, n18207,
         n18208, n18209, n18210, n18211, n18212, n18213, n18214, n18215,
         n18216, n18217, n18218, n18219, n18220, n18221, n18222, n18223,
         n18224, n18225, n18226, n18227, n18228, n18229, n18230, n18231,
         n18232, n18233, n18234, n18235, n18236, n18237, n18238, n18239,
         n18240, n18241, n18242, n18243, n18244, n18245, n18246, n18247,
         n18248, n18249, n18250, n18251, n18252, n18253, n18254, n18255,
         n18256, n18257, n18258, n18259, n18260, n18261, n18262, n18263,
         n18264, n18265, n18266, n18267, n18268, n18269, n18270, n18271,
         n18272, n18273, n18274, n18275, n18276, n18277, n18278, n18279,
         n18280, n18281, n18282, n18283, n18284, n18285, n18286, n18287,
         n18288, n18289, n18290, n18291, n18292, n18293, n18294, n18295,
         n18296, n18297, n18298, n18299, n18300, n18301, n18302, n18303,
         n18304, n18305, n18306, n18307, n18308, n18309, n18310, n18311,
         n18312, n18313, n18314, n18315, n18316, n18317, n18318, n18319,
         n18320, n18321, n18322, n18323, n18324, n18325, n18326, n18327,
         n18328, n18329, n18330, n18331, n18332, n18333, n18334, n18335,
         n18336, n18337, n18338, n18339, n18340, n18341, n18342, n18343,
         n18344, n18345, n18346, n18347, n18348, n18349, n18350, n18351,
         n18352, n18353, n18354, n18355, n18356, n18357, n18358, n18359,
         n18360, n18361, n18362, n18363, n18364, n18365, n18366, n18367,
         n18368, n18369, n18370, n18371, n18372, n18373, n18374, n18375,
         n18376, n18377, n18378, n18379, n18380, n18381, n18382, n18383,
         n18384, n18385, n18386, n18387, n18388, n18389, n18390, n18391,
         n18392, n18393, n18394, n18395, n18396, n18397, n18398, n18399,
         n18400, n18401, n18402, n18403, n18404, n18405, n18406, n18407,
         n18408, n18409, n18410, n18411, n18412, n18413, n18414, n18415,
         n18416, n18417, n18418, n18419, n18420, n18421, n18422, n18423,
         n18424, n18425, n18426, n18427, n18428, n18429, n18430, n18431,
         n18432, n18433, n18434, n18435, n18436, n18437, n18438, n18439,
         n18440, n18441, n18442, n18443, n18444, n18445, n18446, n18447,
         n18448, n18449, n18450, n18451, n18452, n18453, n18454, n18455,
         n18456, n18457, n18458, n18459, n18460, n18461, n18462, n18463,
         n18464, n18465, n18466, n18467, n18468, n18469, n18470, n18471,
         n18472, n18473, n18474, n18475, n18476, n18477, n18478, n18479,
         n18480, n18481, n18482, n18483, n18484, n18485, n18486, n18487,
         n18488, n18489, n18490, n18491, n18492, n18493, n18494, n18495,
         n18496, n18497, n18498, n18499, n18500, n18501, n18502, n18503,
         n18504, n18505, n18506, n18507, n18508, n18509, n18510, n18511,
         n18512, n18513, n18514, n18515, n18516, n18517, n18518, n18519,
         n18520, n18521, n18522, n18523, n18524, n18525, n18526, n18527,
         n18528, n18529, n18530, n18531, n18532, n18533, n18534, n18535,
         n18536, n18537, n18538, n18539, n18540, n18541, n18542, n18543,
         n18544, n18545, n18546, n18547, n18548, n18549, n18550, n18551,
         n18552, n18553, n18554, n18555, n18556, n18557, n18558, n18559,
         n18560, n18561, n18562, n18563, n18564, n18565, n18566, n18567,
         n18568, n18569, n18570, n18571, n18572, n18573, n18574, n18575,
         n18576, n18577, n18578, n18579, n18580, n18581, n18582, n18583,
         n18584, n18585, n18586, n18587, n18588, n18589, n18590, n18591,
         n18592, n18593, n18594, n18595, n18596, n18597, n18598, n18599,
         n18600, n18601, n18602, n18603, n18604, n18605, n18606, n18607,
         n18608, n18609, n18610, n18611, n18612, n18613, n18614, n18615,
         n18616, n18617, n18618, n18619, n18620, n18621, n18622, n18623,
         n18624, n18625, n18626, n18627, n18628, n18629, n18630, n18631,
         n18632, n18633, n18634, n18635, n18636, n18637, n18638, n18639,
         n18640, n18641, n18642, n18643, n18644, n18645, n18646, n18647,
         n18648, n18649, n18650, n18651, n18652, n18653, n18654, n18655,
         n18656, n18657, n18658, n18659, n18660, n18661, n18662, n18663,
         n18664, n18665, n18666, n18667, n18668, n18669, n18670, n18671,
         n18672, n18673, n18674, n18675, n18676, n18677, n18678, n18679,
         n18680, n18681, n18682, n18683, n18684, n18685, n18686, n18687,
         n18688, n18689, n18690, n18691, n18692, n18693, n18694, n18695,
         n18696, n18697, n18698, n18699, n18700, n18701, n18702, n18703,
         n18704, n18705, n18706, n18707, n18708, n18709, n18710, n18711,
         n18712, n18713, n18714, n18715, n18716, n18717, n18718, n18719,
         n18720, n18721, n18722, n18723, n18724, n18725, n18726, n18727,
         n18728, n18729, n18730, n18731, n18732, n18733, n18734, n18735,
         n18736, n18737, n18738, n18739, n18740, n18741, n18742, n18743,
         n18744, n18745, n18746, n18747, n18748, n18749, n18750, n18751,
         n18752, n18753, n18754, n18755, n18756, n18757, n18758, n18759,
         n18760, n18761, n18762, n18763, n18764, n18765, n18766, n18767,
         n18768, n18769, n18770, n18771, n18772, n18773, n18774, n18775,
         n18776, n18777, n18778, n18779, n18780, n18781, n18782, n18783,
         n18784, n18785, n18786, n18787, n18788, n18789, n18790, n18791,
         n18792, n18793, n18794, n18795, n18796, n18797, n18798, n18799,
         n18800, n18801, n18802, n18803, n18804, n18805, n18806, n18807,
         n18808, n18809, n18810, n18811, n18812, n18813, n18814, n18815,
         n18816, n18817, n18818, n18819, n18820, n18821, n18822, n18823,
         n18824, n18825, n18826, n18827, n18828, n18829, n18830, n18831,
         n18832, n18833, n18834, n18835, n18836, n18837, n18838, n18839,
         n18840, n18841, n18842, n18843, n18844, n18845, n18846, n18847,
         n18848, n18849, n18850, n18851, n18852, n18853, n18854, n18855,
         n18856, n18857, n18858, n18859, n18860, n18861, n18862, n18863,
         n18864, n18865, n18866, n18867, n18868, n18869, n18870, n18871,
         n18872, n18873, n18874, n18875, n18876, n18877, n18878, n18879,
         n18880, n18881, n18882, n18883, n18884, n18885, n18886, n18887,
         n18888, n18889, n18890, n18891, n18892, n18893, n18894, n18895,
         n18896, n18897, n18898, n18899, n18900, n18901, n18902, n18903,
         n18904, n18905, n18906, n18907, n18908, n18909, n18910, n18911,
         n18912, n18913, n18914, n18915, n18916, n18917, n18918, n18919,
         n18920, n18921, n18922, n18923, n18924, n18925, n18926, n18927,
         n18928, n18929, n18930, n18931, n18932, n18933, n18934, n18935,
         n18936, n18937, n18938, n18939, n18940, n18941, n18942, n18943,
         n18944, n18945, n18946, n18947, n18948, n18949, n18950, n18951,
         n18952, n18953, n18954, n18955, n18956, n18957, n18958, n18959,
         n18960, n18961, n18962, n18963, n18964, n18965, n18966, n18967,
         n18968, n18969, n18970, n18971, n18972, n18973, n18974, n18975,
         n18976, n18977, n18978, n18979, n18980, n18981, n18982, n18983,
         n18984, n18985, n18986, n18987, n18988, n18989, n18990, n18991,
         n18992, n18993, n18994, n18995, n18996, n18997, n18998, n18999,
         n19000, n19001, n19002, n19003, n19004, n19005, n19006, n19007,
         n19008, n19009, n19010, n19011, n19012, n19013, n19014, n19015,
         n19016, n19017, n19018, n19019, n19020, n19021, n19022, n19023,
         n19024, n19025, n19026, n19027, n19028, n19029, n19030, n19031,
         n19032, n19033, n19034, n19035, n19036, n19037, n19038, n19039,
         n19040, n19041, n19042, n19043, n19044, n19045, n19046, n19047,
         n19048, n19049, n19050, n19051, n19052, n19053, n19054, n19055,
         n19056, n19057, n19058, n19059, n19060, n19061, n19062, n19063,
         n19064, n19065, n19066, n19067, n19068, n19069, n19070, n19071,
         n19072, n19073, n19074, n19075, n19076, n19077, n19078, n19079,
         n19080, n19081, n19082, n19083, n19084, n19085, n19086, n19087,
         n19088, n19089, n19090, n19091, n19092, n19093, n19094, n19095,
         n19096, n19097, n19098, n19099, n19100, n19101, n19102, n19103,
         n19104, n19105, n19106, n19107, n19108, n19109, n19110, n19111,
         n19112, n19113, n19114, n19115, n19116, n19117, n19118, n19119,
         n19120, n19121, n19122, n19123, n19124, n19125, n19126, n19127,
         n19128, n19129, n19130, n19131, n19132, n19133, n19134, n19135,
         n19136, n19137, n19138, n19139, n19140, n19141, n19142, n19143,
         n19144, n19145, n19146, n19147, n19148, n19149, n19150, n19151,
         n19152, n19153, n19154, n19155, n19156, n19157, n19158, n19159,
         n19160, n19161, n19162, n19163, n19164, n19165, n19166, n19167,
         n19168, n19169, n19170, n19171, n19172, n19173, n19174, n19175,
         n19176, n19177, n19178, n19179, n19180, n19181, n19182, n19183,
         n19184, n19185, n19186, n19187, n19188, n19189, n19190, n19191,
         n19192, n19193, n19194, n19195, n19196, n19197, n19198, n19199,
         n19200, n19201, n19202, n19203, n19204, n19205, n19206, n19207,
         n19208, n19209, n19210, n19211, n19212, n19213, n19214, n19215,
         n19216, n19217, n19218, n19219, n19220, n19221, n19222, n19223,
         n19224, n19225, n19226, n19227, n19228, n19229, n19230, n19231,
         n19232, n19233, n19234, n19235, n19236, n19237, n19238, n19239,
         n19240, n19241, n19242, n19243, n19244, n19245, n19246, n19247,
         n19248, n19249, n19250, n19251, n19252, n19253, n19254, n19255,
         n19256, n19257, n19258, n19259, n19260, n19261, n19262, n19263,
         n19264, n19265, n19266, n19267, n19268, n19269, n19270, n19271,
         n19272, n19273, n19274, n19275, n19276, n19277, n19278, n19279,
         n19280, n19281, n19282, n19283, n19284, n19285, n19286, n19287,
         n19288, n19289, n19290, n19291, n19292, n19293, n19294, n19295,
         n19296, n19297, n19298, n19299, n19300, n19301, n19302, n19303,
         n19304, n19305, n19306, n19307, n19308, n19309, n19310, n19311,
         n19312, n19313, n19314, n19315, n19316, n19317, n19318, n19319,
         n19320, n19321, n19322, n19323, n19324, n19325, n19326, n19327,
         n19328, n19329, n19330, n19331, n19332, n19333, n19334, n19335,
         n19336, n19337, n19338, n19339, n19340, n19341, n19342, n19343,
         n19344, n19345, n19346, n19347, n19348, n19349, n19350, n19351,
         n19352, n19353, n19354, n19355, n19356, n19357, n19358, n19359,
         n19360, n19361, n19362, n19363, n19364, n19365, n19366, n19367,
         n19368, n19369, n19370, n19371, n19372, n19373, n19374, n19375,
         n19376, n19377, n19378, n19379, n19380, n19381, n19382, n19383,
         n19384, n19385, n19386, n19387, n19388, n19389, n19390, n19391,
         n19392, n19393, n19394, n19395, n19396, n19397, n19398, n19399,
         n19400, n19401, n19402, n19403, n19404, n19405, n19406, n19407,
         n19408, n19409, n19410, n19411, n19412, n19413, n19414, n19415,
         n19416, n19417, n19418, n19419, n19420, n19421, n19422, n19423,
         n19424, n19425, n19426, n19427, n19428, n19429, n19430, n19431,
         n19432, n19433, n19434, n19435, n19436, n19437, n19438, n19439,
         n19440, n19441, n19442, n19443, n19444, n19445, n19446, n19447,
         n19448, n19449, n19450, n19451, n19452, n19453, n19454, n19455,
         n19456, n19457, n19458, n19459, n19460, n19461, n19462, n19463,
         n19464, n19465, n19466, n19467, n19468, n19469, n19470, n19471,
         n19472, n19473, n19474, n19475, n19476, n19477, n19478, n19479,
         n19480, n19481, n19482, n19483, n19484, n19485, n19486, n19487,
         n19488, n19489, n19490, n19491, n19492, n19493, n19494, n19495,
         n19496, n19497, n19498, n19499, n19500, n19501, n19502, n19503,
         n19504, n19505, n19506, n19507, n19508, n19509, n19510, n19511,
         n19512, n19513, n19514, n19515, n19516, n19517, n19518, n19519,
         n19520, n19521, n19522, n19523, n19524, n19525, n19526, n19527,
         n19528, n19529, n19530, n19531, n19532, n19533, n19534, n19535,
         n19536, n19537, n19538, n19539, n19540, n19541, n19542, n19543,
         n19544, n19545, n19546, n19547, n19548, n19549, n19550, n19551,
         n19552, n19553, n19554, n19555, n19556, n19557, n19558, n19559,
         n19560, n19561, n19562, n19563, n19564, n19565, n19566, n19567,
         n19568, n19569, n19570, n19571, n19572, n19573, n19574, n19575,
         n19576, n19577, n19578, n19579, n19580, n19581, n19582, n19583,
         n19584, n19585, n19586, n19587, n19588, n19589, n19590, n19591,
         n19592, n19593, n19594, n19595, n19596, n19597, n19598, n19599,
         n19600, n19601, n19602, n19603, n19604, n19605, n19606, n19607,
         n19608, n19609, n19610, n19611, n19612, n19613, n19614, n19615,
         n19616, n19617, n19618, n19619, n19620, n19621, n19622, n19623,
         n19624, n19625, n19626, n19627, n19628, n19629, n19630, n19631,
         n19632, n19633, n19634, n19635, n19636, n19637, n19638, n19639,
         n19640, n19641, n19642, n19643, n19644, n19645, n19646, n19647,
         n19648, n19649, n19650, n19651, n19652, n19653, n19654, n19655,
         n19656, n19657, n19658, n19659, n19660, n19661, n19662, n19663,
         n19664, n19665, n19666, n19667, n19668, n19669, n19670, n19671,
         n19672, n19673, n19674, n19675, n19676, n19677, n19678, n19679,
         n19680, n19681, n19682, n19683, n19684, n19685, n19686, n19687,
         n19688, n19689, n19690, n19691, n19692, n19693, n19694, n19695,
         n19696, n19697, n19698, n19699, n19700, n19701, n19702, n19703,
         n19704, n19705, n19706, n19707, n19708, n19709, n19710, n19711,
         n19712, n19713, n19714, n19715, n19716, n19717, n19718, n19719,
         n19720, n19721, n19722, n19723, n19724, n19725, n19726, n19727,
         n19728, n19729, n19730, n19731, n19732, n19733, n19734, n19735,
         n19736, n19737, n19738, n19739, n19740, n19741, n19742, n19743,
         n19744, n19745, n19746, n19747, n19748, n19749, n19750, n19751,
         n19752, n19753, n19754, n19755, n19756, n19757, n19758, n19759,
         n19760, n19761, n19762, n19763, n19764, n19765, n19766, n19767,
         n19768, n19769, n19770, n19771, n19772, n19773, n19774, n19775,
         n19776, n19777, n19778, n19779, n19780, n19781, n19782, n19783,
         n19784, n19785, n19786, n19787, n19788, n19789, n19790, n19791,
         n19792, n19793, n19794, n19795, n19796, n19797, n19798, n19799,
         n19800, n19801, n19802, n19803, n19804, n19805, n19806, n19807,
         n19808, n19809, n19810, n19811, n19812, n19813, n19814, n19815,
         n19816, n19817, n19818, n19819, n19820, n19821, n19822, n19823,
         n19824, n19825, n19826, n19827, n19828, n19829, n19830, n19831,
         n19832, n19833, n19834, n19835, n19836, n19837, n19838, n19839,
         n19840, n19841, n19842, n19843, n19844, n19845, n19846, n19847,
         n19848, n19849, n19850, n19851, n19852, n19853, n19854, n19855,
         n19856, n19857, n19858, n19859, n19860, n19861, n19862, n19863,
         n19864, n19865, n19866, n19867, n19868, n19869, n19870, n19871,
         n19872, n19873, n19874, n19875, n19876, n19877, n19878, n19879,
         n19880, n19881, n19882, n19883, n19884, n19885, n19886, n19887,
         n19888, n19889, n19890, n19891, n19892, n19893, n19894, n19895,
         n19896, n19897, n19898, n19899, n19900, n19901, n19902, n19903,
         n19904, n19905, n19906, n19907, n19908, n19909, n19910, n19911,
         n19912, n19913, n19914, n19915, n19916, n19917, n19918, n19919,
         n19920, n19921, n19922, n19923, n19924, n19925, n19926, n19927,
         n19928, n19929, n19930, n19931, n19932, n19933, n19934, n19935,
         n19936, n19937, n19938, n19939, n19940, n19941, n19942, n19943,
         n19944, n19945, n19946, n19947, n19948, n19949, n19950, n19951,
         n19952, n19953, n19954, n19955, n19956, n19957, n19958, n19959,
         n19960, n19961, n19962, n19963, n19964, n19965, n19966, n19967,
         n19968, n19969, n19970, n19971, n19972, n19973, n19974, n19975,
         n19976, n19977, n19978, n19979, n19980, n19981, n19982, n19983,
         n19984, n19985, n19986, n19987, n19988, n19989, n19990, n19991,
         n19992, n19993, n19994, n19995, n19996, n19997, n19998, n19999,
         n20000, n20001, n20002, n20003, n20004, n20005, n20006, n20007,
         n20008, n20009, n20010, n20011, n20012, n20013, n20014, n20015,
         n20016, n20017, n20018, n20019, n20020, n20021, n20022, n20023,
         n20024, n20025, n20026, n20027, n20028, n20029, n20030, n20031,
         n20032, n20033, n20034, n20035, n20036, n20037, n20038, n20039,
         n20040, n20041, n20042, n20043, n20044, n20045, n20046, n20047,
         n20048, n20049, n20050, n20051, n20052, n20053, n20054, n20055,
         n20056, n20057, n20058, n20059, n20060, n20061, n20062, n20063,
         n20064, n20065, n20066, n20067, n20068, n20069, n20070, n20071,
         n20072, n20073, n20074, n20075, n20076, n20077, n20078, n20079,
         n20080, n20081, n20082, n20083, n20084, n20085, n20086, n20087,
         n20088, n20089, n20090, n20091, n20092, n20093, n20094, n20095,
         n20096, n20097, n20098, n20099, n20100, n20101, n20102, n20103,
         n20104, n20105, n20106, n20107, n20108, n20109, n20110, n20111,
         n20112, n20113, n20114, n20115, n20116, n20117, n20118, n20119,
         n20120, n20121, n20122, n20123, n20124, n20125, n20126, n20127,
         n20128, n20129, n20130, n20131, n20132, n20133, n20134, n20135,
         n20136, n20137, n20138, n20139, n20140, n20141, n20142, n20143,
         n20144, n20145, n20146, n20147, n20148, n20149, n20150, n20151,
         n20152, n20153, n20154, n20155, n20156, n20157, n20158, n20159,
         n20160, n20161, n20162, n20163, n20164, n20165, n20166, n20167,
         n20168, n20169, n20170, n20171, n20172, n20173, n20174, n20175,
         n20176, n20177, n20178, n20179, n20180, n20181, n20182, n20183,
         n20184, n20185, n20186, n20187, n20188, n20189, n20190, n20191,
         n20192, n20193, n20194, n20195, n20196, n20197, n20198, n20199,
         n20200, n20201, n20202, n20203, n20204, n20205, n20206, n20207,
         n20208, n20209, n20210, n20211, n20212, n20213, n20214, n20215,
         n20216, n20217, n20218, n20219, n20220, n20221, n20222, n20223,
         n20224, n20225, n20226, n20227, n20228, n20229, n20230, n20231,
         n20232, n20233, n20234, n20235, n20236, n20237, n20238, n20239,
         n20240, n20241, n20242, n20243, n20244, n20245, n20246, n20247,
         n20248, n20249, n20250, n20251, n20252, n20253, n20254, n20255,
         n20256, n20257, n20258, n20259, n20260, n20261, n20262, n20263,
         n20264, n20265, n20266, n20267, n20268, n20269, n20270, n20271,
         n20272, n20273, n20274, n20275, n20276, n20277, n20278, n20279,
         n20280, n20281, n20282, n20283, n20284, n20285, n20286, n20287,
         n20288, n20289, n20290, n20291, n20292, n20293, n20294, n20295,
         n20296, n20297, n20298, n20299, n20300, n20301, n20302, n20303,
         n20304, n20305, n20306, n20307, n20308, n20309, n20310, n20311,
         n20312, n20313, n20314, n20315, n20316, n20317, n20318, n20319,
         n20320, n20321, n20322, n20323, n20324, n20325, n20326, n20327,
         n20328, n20329, n20330, n20331, n20332, n20333, n20334, n20335,
         n20336, n20337, n20338, n20339, n20340, n20341, n20342, n20343,
         n20344, n20345, n20346, n20347, n20348, n20349, n20350, n20351,
         n20352, n20353, n20354, n20355, n20356, n20357, n20358, n20359,
         n20360, n20361, n20362, n20363, n20364, n20365, n20366, n20367,
         n20368, n20369, n20370, n20371, n20372, n20373, n20374, n20375,
         n20376, n20377, n20378, n20379, n20380, n20381, n20382, n20383,
         n20384, n20385, n20386, n20387, n20388, n20389, n20390, n20391,
         n20392, n20393, n20394, n20395, n20396, n20397, n20398, n20399,
         n20400, n20401, n20402, n20403, n20404, n20405, n20406, n20407,
         n20408, n20409, n20410, n20411, n20412, n20413, n20414, n20415,
         n20416, n20417, n20418, n20419, n20420, n20421, n20422, n20423,
         n20424, n20425, n20426, n20427, n20428, n20429, n20430, n20431,
         n20432, n20433, n20434, n20435, n20436, n20437, n20438, n20439,
         n20440, n20441, n20442, n20443, n20444, n20445, n20446, n20447,
         n20448, n20449, n20450, n20451, n20452, n20453, n20454, n20455,
         n20456, n20457, n20458, n20459, n20460, n20461, n20462, n20463,
         n20464, n20465, n20466, n20467, n20468, n20469, n20470, n20471,
         n20472, n20473, n20474, n20475, n20476, n20477, n20478, n20479,
         n20480, n20481, n20482, n20483, n20484, n20485, n20486, n20487,
         n20488, n20489, n20490, n20491, n20492, n20493, n20494, n20495,
         n20496, n20497, n20498, n20499, n20500, n20501, n20502, n20503,
         n20504, n20505, n20506, n20507, n20508, n20509, n20510, n20511,
         n20512, n20513, n20514, n20515, n20516, n20517, n20518, n20519,
         n20520, n20521, n20522, n20523, n20524, n20525, n20526, n20527,
         n20528, n20529, n20530, n20531, n20532, n20533, n20534, n20535,
         n20536, n20537, n20538, n20539, n20540, n20541, n20542, n20543,
         n20544, n20545, n20546, n20547, n20548, n20549, n20550, n20551,
         n20552, n20553, n20554, n20555, n20556, n20557, n20558, n20559,
         n20560, n20561, n20562, n20563, n20564, n20565, n20566, n20567,
         n20568, n20569, n20570, n20571, n20572, n20573, n20574, n20575,
         n20576, n20577, n20578, n20579, n20580, n20581, n20582, n20583,
         n20584, n20585, n20586, n20587, n20588, n20589, n20590, n20591,
         n20592, n20593, n20594, n20595, n20596, n20597, n20598, n20599,
         n20600, n20601, n20602, n20603, n20604, n20605, n20606, n20607,
         n20608, n20609, n20610, n20611, n20612, n20613, n20614, n20615,
         n20616, n20617, n20618, n20619, n20620, n20621, n20622, n20623,
         n20624, n20625, n20626, n20627, n20628, n20629, n20630, n20631,
         n20632, n20633, n20634, n20635, n20636, n20637, n20638, n20639,
         n20640, n20641, n20642, n20643, n20644, n20645, n20646, n20647,
         n20648, n20649, n20650, n20651, n20652, n20653, n20654, n20655,
         n20656, n20657, n20658, n20659, n20660, n20661, n20662, n20663,
         n20664, n20665, n20666, n20667, n20668, n20669, n20670, n20671,
         n20672, n20673, n20674, n20675, n20676, n20677, n20678, n20679,
         n20680, n20681, n20682, n20683, n20684, n20685, n20686, n20687,
         n20688, n20689, n20690, n20691, n20692, n20693, n20694, n20695,
         n20696, n20697, n20698, n20699, n20700, n20701, n20702, n20703,
         n20704, n20705, n20706, n20707, n20708, n20709, n20710, n20711,
         n20712, n20713, n20714, n20715, n20716, n20717, n20718, n20719,
         n20720, n20721, n20722, n20723, n20724, n20725, n20726, n20727,
         n20728, n20729, n20730, n20731, n20732, n20733, n20734, n20735,
         n20736, n20737, n20738, n20739, n20740, n20741, n20742, n20743,
         n20744, n20745, n20746, n20747, n20748, n20749, n20750, n20751,
         n20752, n20753, n20754, n20755, n20756, n20757, n20758, n20759,
         n20760, n20761, n20762, n20763, n20764, n20765, n20766, n20767,
         n20768, n20769, n20770, n20771, n20772, n20773, n20774, n20775,
         n20776, n20777, n20778, n20779, n20780, n20781, n20782, n20783,
         n20784, n20785, n20786, n20787, n20788, n20789, n20790, n20791,
         n20792, n20793, n20794, n20795, n20796, n20797, n20798, n20799,
         n20800, n20801, n20802, n20803, n20804, n20805, n20806, n20807,
         n20808, n20809, n20810, n20811, n20812, n20813, n20814, n20815,
         n20816, n20817, n20818, n20819, n20820, n20821, n20822, n20823,
         n20824, n20825, n20826, n20827, n20828, n20829, n20830, n20831,
         n20832, n20833, n20834, n20835, n20836, n20837, n20838, n20839,
         n20840, n20841, n20842, n20843, n20844, n20845, n20846, n20847,
         n20848, n20849, n20850, n20851, n20852, n20853, n20854, n20855,
         n20856, n20857, n20858, n20859, n20860, n20861, n20862, n20863,
         n20864, n20865, n20866, n20867, n20868, n20869, n20870, n20871,
         n20872, n20873, n20874, n20875, n20876, n20877, n20878, n20879,
         n20880, n20881, n20882, n20883, n20884, n20885, n20886, n20887,
         n20888, n20889, n20890, n20891, n20892, n20893, n20894, n20895,
         n20896, n20897, n20898, n20899, n20900, n20901, n20902, n20903,
         n20904, n20905, n20906, n20907, n20908, n20909, n20910, n20911,
         n20912, n20913, n20914, n20915, n20916, n20917, n20918, n20919,
         n20920, n20921, n20922, n20923, n20924, n20925, n20926, n20927,
         n20928, n20929, n20930, n20931, n20932, n20933, n20934, n20935,
         n20936, n20937, n20938, n20939, n20940, n20941, n20942, n20943,
         n20944, n20945, n20946, n20947, n20948, n20949, n20950, n20951,
         n20952, n20953, n20954, n20955, n20956, n20957, n20958, n20959,
         n20960, n20961, n20962, n20963, n20964, n20965, n20966, n20967,
         n20968, n20969, n20970, n20971, n20972, n20973, n20974, n20975,
         n20976, n20977, n20978, n20979, n20980, n20981, n20982, n20983,
         n20984, n20985, n20986, n20987, n20988, n20989, n20990, n20991,
         n20992, n20993, n20994, n20995, n20996, n20997, n20998, n20999,
         n21000, n21001, n21002, n21003, n21004, n21005, n21006, n21007,
         n21008, n21009, n21010, n21011, n21012, n21013, n21014, n21015,
         n21016, n21017, n21018, n21019, n21020, n21021, n21022, n21023,
         n21024, n21025, n21026, n21027, n21028, n21029, n21030, n21031,
         n21032, n21033, n21034, n21035, n21036, n21037, n21038, n21039,
         n21040, n21041, n21042, n21043, n21044, n21045, n21046, n21047,
         n21048, n21049, n21050, n21051, n21052, n21053, n21054, n21055,
         n21056, n21057, n21058, n21059, n21060, n21061, n21062, n21063,
         n21064, n21065, n21066, n21067, n21068, n21069, n21070, n21071,
         n21072, n21073, n21074, n21075, n21076, n21077, n21078, n21079,
         n21080, n21081, n21082, n21083, n21084, n21085, n21086, n21087,
         n21088, n21089, n21090, n21091, n21092, n21093, n21094, n21095,
         n21096, n21097, n21098, n21099, n21100, n21101, n21102, n21103,
         n21104, n21105, n21106, n21107, n21108, n21109, n21110, n21111,
         n21112, n21113, n21114, n21115, n21116, n21117, n21118, n21119,
         n21120, n21121, n21122, n21123, n21124, n21125, n21126, n21127,
         n21128, n21129, n21130, n21131, n21132, n21133, n21134, n21135,
         n21136, n21137, n21138, n21139, n21140, n21141, n21142, n21143,
         n21144, n21145, n21146, n21147, n21148, n21149, n21150, n21151,
         n21152, n21153, n21154, n21155, n21156, n21157, n21158, n21159,
         n21160, n21161, n21162, n21163, n21164, n21165, n21166, n21167,
         n21168, n21169, n21170, n21171, n21172, n21173, n21174, n21175,
         n21176, n21177, n21178, n21179, n21180, n21181, n21182, n21183,
         n21184, n21185, n21186, n21187, n21188, n21189, n21190, n21191,
         n21192, n21193, n21194, n21195, n21196, n21197, n21198, n21199,
         n21200, n21201, n21202, n21203, n21204, n21205, n21206, n21207,
         n21208, n21209, n21210, n21211, n21212, n21213, n21214, n21215,
         n21216, n21217, n21218, n21219, n21220, n21221, n21222, n21223,
         n21224, n21225, n21226, n21227, n21228, n21229, n21230, n21231,
         n21232, n21233, n21234, n21235, n21236, n21237, n21238, n21239,
         n21240, n21241, n21242, n21243, n21244, n21245, n21246, n21247,
         n21248, n21249, n21250, n21251, n21252, n21253, n21254, n21255,
         n21256, n21257, n21258, n21259, n21260, n21261, n21262, n21263,
         n21264, n21265, n21266, n21267, n21268, n21269, n21270, n21271,
         n21272, n21273, n21274, n21275, n21276, n21277, n21278, n21279,
         n21280, n21281, n21282, n21283, n21284, n21285, n21286, n21287,
         n21288, n21289, n21290, n21291, n21292, n21293, n21294, n21295,
         n21296, n21297, n21298, n21299, n21300, n21301, n21302, n21303,
         n21304, n21305, n21306, n21307, n21308, n21309, n21310, n21311,
         n21312, n21313, n21314, n21315, n21316, n21317, n21318, n21319,
         n21320, n21321, n21322, n21323, n21324, n21325, n21326, n21327,
         n21328, n21329, n21330, n21331, n21332, n21333, n21334, n21335,
         n21336, n21337, n21338, n21339, n21340, n21341, n21342, n21343,
         n21344, n21345, n21346, n21347, n21348, n21349, n21350, n21351,
         n21352, n21353, n21354, n21355, n21356, n21357, n21358, n21359,
         n21360, n21361, n21362, n21363, n21364, n21365, n21366, n21367,
         n21368, n21369, n21370, n21371, n21372, n21373, n21374, n21375,
         n21376, n21377, n21378, n21379, n21380, n21381, n21382, n21383,
         n21384, n21385, n21386, n21387, n21388, n21389, n21390, n21391,
         n21392, n21393, n21394, n21395, n21396, n21397, n21398, n21399,
         n21400, n21401, n21402, n21403, n21404, n21405, n21406, n21407,
         n21408, n21409, n21410, n21411, n21412, n21413, n21414, n21415,
         n21416, n21417, n21418, n21419, n21420, n21421, n21422, n21423,
         n21424, n21425, n21426, n21427, n21428, n21429, n21430, n21431,
         n21432, n21433, n21434, n21435, n21436, n21437, n21438, n21439,
         n21440, n21441, n21442, n21443, n21444, n21445, n21446, n21447,
         n21448, n21449, n21450, n21451, n21452, n21453, n21454, n21455,
         n21456, n21457, n21458, n21459, n21460, n21461, n21462, n21463,
         n21464, n21465, n21466, n21467, n21468, n21469, n21470, n21471,
         n21472, n21473, n21474, n21475, n21476, n21477, n21478, n21479,
         n21480, n21481, n21482, n21483, n21484, n21485, n21486, n21487,
         n21488, n21489, n21490, n21491, n21492, n21493, n21494, n21495,
         n21496, n21497, n21498, n21499, n21500, n21501, n21502, n21503,
         n21504, n21505, n21506, n21507, n21508, n21509, n21510, n21511,
         n21512, n21513, n21514, n21515, n21516, n21517, n21518, n21519,
         n21520, n21521, n21522, n21523, n21524, n21525, n21526, n21527,
         n21528, n21529, n21530, n21531, n21532, n21533, n21534, n21535,
         n21536, n21537, n21538, n21539, n21540, n21541, n21542, n21543,
         n21544, n21545, n21546, n21547, n21548, n21549, n21550, n21551,
         n21552, n21553, n21554, n21555, n21556, n21557, n21558, n21559,
         n21560, n21561, n21562, n21563, n21564, n21565, n21566, n21567,
         n21568, n21569, n21570, n21571, n21572, n21573, n21574, n21575,
         n21576, n21577, n21578, n21579, n21580, n21581, n21582, n21583,
         n21584, n21585, n21586, n21587, n21588, n21589, n21590, n21591,
         n21592, n21593, n21594, n21595, n21596, n21597, n21598, n21599,
         n21600, n21601, n21602, n21603, n21604, n21605, n21606, n21607,
         n21608, n21609, n21610, n21611, n21612, n21613, n21614, n21615,
         n21616, n21617, n21618, n21619, n21620, n21621, n21622, n21623,
         n21624, n21625, n21626, n21627, n21628, n21629, n21630, n21631,
         n21632, n21633, n21634, n21635, n21636, n21637, n21638, n21639,
         n21640, n21641, n21642, n21643, n21644, n21645, n21646, n21647,
         n21648, n21649, n21650, n21651, n21652, n21653, n21654, n21655,
         n21656, n21657, n21658, n21659, n21660, n21661, n21662, n21663,
         n21664, n21665, n21666, n21667, n21668, n21669, n21670, n21671,
         n21672, n21673, n21674, n21675, n21676, n21677, n21678, n21679,
         n21680, n21681, n21682, n21683, n21684, n21685, n21686, n21687,
         n21688, n21689, n21690, n21691, n21692, n21693, n21694, n21695,
         n21696, n21697, n21698, n21699, n21700, n21701, n21702, n21703,
         n21704, n21705, n21706, n21707, n21708, n21709, n21710, n21711,
         n21712, n21713, n21714, n21715, n21716, n21717, n21718, n21719,
         n21720, n21721, n21722, n21723, n21724, n21725, n21726, n21727,
         n21728, n21729, n21730, n21731, n21732, n21733, n21734, n21735,
         n21736, n21737, n21738, n21739, n21740, n21741, n21742, n21743,
         n21744, n21745, n21746, n21747, n21748, n21749, n21750, n21751,
         n21752, n21753, n21754, n21755, n21756, n21757, n21758, n21759,
         n21760, n21761, n21762, n21763, n21764, n21765, n21766, n21767,
         n21768, n21769, n21770, n21771, n21772, n21773, n21774, n21775,
         n21776, n21777, n21778, n21779, n21780, n21781, n21782, n21783,
         n21784, n21785, n21786, n21787, n21788, n21789, n21790, n21791,
         n21792, n21793, n21794, n21795, n21796, n21797, n21798, n21799,
         n21800, n21801, n21802, n21803, n21804, n21805, n21806, n21807,
         n21808, n21809, n21810, n21811, n21812, n21813, n21814, n21815,
         n21816, n21817, n21818, n21819, n21820, n21821, n21822, n21823,
         n21824, n21825, n21826, n21827, n21828, n21829, n21830, n21831,
         n21832, n21833, n21834, n21835, n21836, n21837, n21838, n21839,
         n21840, n21841, n21842, n21843, n21844, n21845, n21846, n21847,
         n21848, n21849, n21850, n21851, n21852, n21853, n21854, n21855,
         n21856, n21857, n21858, n21859, n21860, n21861, n21862, n21863,
         n21864, n21865, n21866, n21867, n21868, n21869, n21870, n21871,
         n21872, n21873, n21874, n21875, n21876, n21877, n21878, n21879,
         n21880, n21881, n21882, n21883, n21884, n21885, n21886, n21887,
         n21888, n21889, n21890, n21891, n21892, n21893, n21894, n21895,
         n21896, n21897, n21898, n21899, n21900, n21901, n21902, n21903,
         n21904, n21905, n21906, n21907, n21908, n21909, n21910, n21911,
         n21912, n21913, n21914, n21915, n21916, n21917, n21918, n21919,
         n21920, n21921, n21922, n21923, n21924, n21925, n21926, n21927,
         n21928, n21929, n21930, n21931, n21932, n21933, n21934, n21935,
         n21936, n21937, n21938, n21939, n21940, n21941, n21942, n21943,
         n21944, n21945, n21946, n21947, n21948, n21949, n21950, n21951,
         n21952, n21953, n21954, n21955, n21956, n21957, n21958, n21959,
         n21960, n21961, n21962, n21963, n21964, n21965, n21966, n21967,
         n21968, n21969, n21970, n21971, n21972, n21973, n21974, n21975,
         n21976, n21977, n21978, n21979, n21980, n21981, n21982, n21983,
         n21984, n21985, n21986, n21987, n21988, n21989, n21990, n21991,
         n21992, n21993, n21994, n21995, n21996, n21997, n21998, n21999,
         n22000, n22001, n22002, n22003, n22004, n22005, n22006, n22007,
         n22008, n22009, n22010, n22011, n22012, n22013, n22014, n22015,
         n22016, n22017, n22018, n22019, n22020, n22021, n22022, n22023,
         n22024, n22025, n22026, n22027, n22028, n22029, n22030, n22031,
         n22032, n22033, n22034, n22035, n22036, n22037, n22038, n22039,
         n22040, n22041, n22042, n22043, n22044, n22045, n22046, n22047,
         n22048, n22049, n22050, n22051, n22052, n22053, n22054, n22055,
         n22056, n22057, n22058, n22059, n22060, n22061, n22062, n22063,
         n22064, n22065, n22066, n22067, n22068, n22069, n22070, n22071,
         n22072, n22073, n22074, n22075, n22076, n22077, n22078, n22079,
         n22080, n22081, n22082, n22083, n22084, n22085, n22086, n22087,
         n22088, n22089, n22090, n22091, n22092, n22093, n22094, n22095,
         n22096, n22097, n22098, n22099, n22100, n22101, n22102, n22103,
         n22104, n22105, n22106, n22107, n22108, n22109, n22110, n22111,
         n22112, n22113, n22114, n22115, n22116, n22117, n22118, n22119,
         n22120, n22121, n22122, n22123, n22124, n22125, n22126, n22127,
         n22128, n22129, n22130, n22131, n22132, n22133, n22134, n22135,
         n22136, n22137, n22138, n22139, n22140, n22141, n22142, n22143,
         n22144, n22145, n22146, n22147, n22148, n22149, n22150, n22151,
         n22152, n22153, n22154, n22155, n22156, n22157, n22158, n22159,
         n22160, n22161, n22162, n22163, n22164, n22165, n22166, n22167,
         n22168, n22169, n22170, n22171, n22172, n22173, n22174, n22175,
         n22176, n22177, n22178, n22179, n22180, n22181, n22182, n22183,
         n22184, n22185, n22186, n22187, n22188, n22189, n22190, n22191,
         n22192, n22193, n22194, n22195, n22196, n22197, n22198, n22199,
         n22200, n22201, n22202, n22203, n22204, n22205, n22206, n22207,
         n22208, n22209, n22210, n22211, n22212, n22213, n22214, n22215,
         n22216, n22217, n22218, n22219, n22220, n22221, n22222, n22223,
         n22224, n22225, n22226, n22227, n22228, n22229, n22230, n22231,
         n22232, n22233, n22234, n22235, n22236, n22237, n22238, n22239,
         n22240, n22241, n22242, n22243, n22244, n22245, n22246, n22247,
         n22248, n22249, n22250, n22251, n22252, n22253, n22254, n22255,
         n22256, n22257, n22258, n22259, n22260, n22261, n22262, n22263,
         n22264, n22265, n22266, n22267, n22268, n22269, n22270, n22271,
         n22272, n22273, n22274, n22275, n22276, n22277, n22278, n22279,
         n22280, n22281, n22282, n22283, n22284, n22285, n22286, n22287,
         n22288, n22289, n22290, n22291, n22292, n22293, n22294, n22295,
         n22296, n22297, n22298, n22299, n22300, n22301, n22302, n22303,
         n22304, n22305, n22306, n22307, n22308, n22309, n22310, n22311,
         n22312, n22313, n22314, n22315, n22316, n22317, n22318, n22319,
         n22320, n22321, n22322, n22323, n22324, n22325, n22326, n22327,
         n22328, n22329, n22330, n22331, n22332, n22333, n22334, n22335,
         n22336, n22337, n22338, n22339, n22340, n22341, n22342, n22343,
         n22344, n22345, n22346, n22347, n22348, n22349, n22350, n22351,
         n22352, n22353, n22354, n22355, n22356, n22357, n22358, n22359,
         n22360, n22361, n22362, n22363, n22364, n22365, n22366, n22367,
         n22368, n22369, n22370, n22371, n22372, n22373, n22374, n22375,
         n22376, n22377, n22378, n22379, n22380, n22381, n22382, n22383,
         n22384, n22385, n22386, n22387, n22388, n22389, n22390, n22391,
         n22392, n22393, n22394, n22395, n22396, n22397, n22398, n22399,
         n22400, n22401, n22402, n22403, n22404, n22405, n22406, n22407,
         n22408, n22409, n22410, n22411, n22412, n22413, n22414, n22415,
         n22416, n22417, n22418, n22419, n22420, n22421, n22422, n22423,
         n22424, n22425, n22426, n22427, n22428, n22429, n22430, n22431,
         n22432, n22433, n22434, n22435, n22436, n22437, n22438, n22439,
         n22440, n22441, n22442, n22443, n22444, n22445, n22446, n22447,
         n22448, n22449, n22450, n22451, n22452, n22453, n22454, n22455,
         n22456, n22457, n22458, n22459, n22460, n22461, n22462, n22463,
         n22464, n22465, n22466, n22467, n22468, n22469, n22470, n22471,
         n22472, n22473, n22474, n22475, n22476, n22477, n22478, n22479,
         n22480, n22481, n22482, n22483, n22484, n22485, n22486, n22487,
         n22488, n22489, n22490, n22491, n22492, n22493, n22494, n22495,
         n22496, n22497, n22498, n22499, n22500, n22501, n22502, n22503,
         n22504, n22505, n22506, n22507, n22508, n22509, n22510, n22511,
         n22512, n22513, n22514, n22515, n22516, n22517, n22518, n22519,
         n22520, n22521, n22522, n22523, n22524, n22525, n22526, n22527,
         n22528, n22529, n22530, n22531, n22532, n22533, n22534, n22535,
         n22536, n22537, n22538, n22539, n22540, n22541, n22542, n22543,
         n22544, n22545, n22546, n22547, n22548, n22549, n22550, n22551,
         n22552, n22553, n22554, n22555, n22556, n22557, n22558, n22559,
         n22560, n22561, n22562, n22563, n22564, n22565, n22566, n22567,
         n22568, n22569, n22570, n22571, n22572, n22573, n22574, n22575,
         n22576, n22577, n22578, n22579, n22580, n22581, n22582, n22583,
         n22584, n22585, n22586, n22587, n22588, n22589, n22590, n22591,
         n22592, n22593, n22594, n22595, n22596, n22597, n22598, n22599,
         n22600, n22601, n22602, n22603, n22604, n22605, n22606, n22607,
         n22608, n22609, n22610, n22611, n22612, n22613, n22614, n22615,
         n22616, n22617, n22618, n22619, n22620, n22621, n22622, n22623,
         n22624, n22625, n22626, n22627, n22628, n22629, n22630, n22631,
         n22632, n22633, n22634, n22635, n22636, n22637, n22638, n22639,
         n22640, n22641, n22642, n22643, n22644, n22645, n22646, n22647,
         n22648, n22649, n22650, n22651, n22652, n22653, n22654, n22655,
         n22656, n22657, n22658, n22659, n22660, n22661, n22662, n22663,
         n22664, n22665, n22666, n22667, n22668, n22669, n22670, n22671,
         n22672, n22673, n22674, n22675, n22676, n22677, n22678, n22679,
         n22680, n22681, n22682, n22683, n22684, n22685, n22686, n22687,
         n22688, n22689, n22690, n22691, n22692, n22693, n22694, n22695,
         n22696, n22697, n22698, n22699, n22700, n22701, n22702, n22703,
         n22704, n22705, n22706, n22707, n22708, n22709, n22710, n22711,
         n22712, n22713, n22714, n22715, n22716, n22717, n22718, n22719,
         n22720, n22721, n22722, n22723, n22724, n22725, n22726, n22727,
         n22728, n22729, n22730, n22731, n22732, n22733, n22734, n22735,
         n22736, n22737, n22738, n22739, n22740, n22741, n22742, n22743,
         n22744, n22745, n22746, n22747, n22748, n22749, n22750, n22751,
         n22752, n22753, n22754, n22755, n22756, n22757, n22758, n22759,
         n22760, n22761, n22762, n22763, n22764, n22765, n22766, n22767,
         n22768, n22769, n22770, n22771, n22772, n22773, n22774, n22775,
         n22776, n22777, n22778, n22779, n22780, n22781, n22782, n22783,
         n22784, n22785, n22786, n22787, n22788, n22789, n22790, n22791,
         n22792, n22793, n22794, n22795, n22796, n22797, n22798, n22799,
         n22800, n22801, n22802, n22803, n22804, n22805, n22806, n22807,
         n22808, n22809, n22810, n22811, n22812, n22813, n22814, n22815,
         n22816, n22817, n22818, n22819, n22820, n22821, n22822, n22823,
         n22824, n22825, n22826, n22827, n22828, n22829, n22830, n22831,
         n22832, n22833, n22834, n22835, n22836, n22837, n22838, n22839,
         n22840, n22841, n22842, n22843, n22844, n22845, n22846, n22847,
         n22848, n22849, n22850, n22851, n22852, n22853, n22854, n22855,
         n22856, n22857, n22858, n22859, n22860, n22861, n22862, n22863,
         n22864, n22865, n22866, n22867, n22868, n22869, n22870, n22871,
         n22872, n22873, n22874, n22875, n22876, n22877, n22878, n22879,
         n22880, n22881, n22882, n22883, n22884, n22885, n22886, n22887,
         n22888, n22889, n22890, n22891, n22892, n22893, n22894, n22895,
         n22896, n22897, n22898, n22899, n22900, n22901, n22902, n22903,
         n22904, n22905, n22906, n22907, n22908, n22909, n22910, n22911,
         n22912, n22913, n22914, n22915, n22916, n22917, n22918, n22919,
         n22920, n22921, n22922, n22923, n22924, n22925, n22926, n22927,
         n22928, n22929, n22930, n22931, n22932, n22933, n22934, n22935,
         n22936, n22937, n22938, n22939, n22940, n22941, n22942, n22943,
         n22944, n22945, n22946, n22947, n22948, n22949, n22950, n22951,
         n22952, n22953, n22954, n22955, n22956, n22957, n22958, n22959,
         n22960, n22961, n22962, n22963, n22964, n22965, n22966, n22967,
         n22968, n22969, n22970, n22971, n22972, n22973, n22974, n22975,
         n22976, n22977, n22978, n22979, n22980, n22981, n22982, n22983,
         n22984, n22985, n22986, n22987, n22988, n22989, n22990, n22991,
         n22992, n22993, n22994, n22995, n22996, n22997, n22998, n22999,
         n23000, n23001, n23002, n23003, n23004, n23005, n23006, n23007,
         n23008, n23009, n23010, n23011, n23012, n23013, n23014, n23015,
         n23016, n23017, n23018, n23019, n23020, n23021, n23022, n23023,
         n23024, n23025, n23026, n23027, n23028, n23029, n23030, n23031,
         n23032, n23033, n23034, n23035, n23036, n23037, n23038, n23039,
         n23040, n23041, n23042, n23043, n23044, n23045, n23046, n23047,
         n23048, n23049, n23050, n23051, n23052, n23053, n23054, n23055,
         n23056, n23057, n23058, n23059, n23060, n23061, n23062, n23063,
         n23064, n23065, n23066, n23067, n23068, n23069, n23070, n23071,
         n23072, n23073, n23074, n23075, n23076, n23077, n23078, n23079,
         n23080, n23081, n23082, n23083, n23084, n23085, n23086, n23087,
         n23088, n23089, n23090, n23091, n23092, n23093, n23094, n23095,
         n23096, n23097, n23098, n23099, n23100, n23101, n23102, n23103,
         n23104, n23105, n23106, n23107, n23108, n23109, n23110, n23111,
         n23112, n23113, n23114, n23115, n23116, n23117, n23118, n23119,
         n23120, n23121, n23122, n23123, n23124, n23125, n23126, n23127,
         n23128, n23129, n23130, n23131, n23132, n23133, n23134, n23135,
         n23136, n23137, n23138, n23139, n23140, n23141, n23142, n23143,
         n23144, n23145, n23146, n23147, n23148, n23149, n23150, n23151,
         n23152, n23153, n23154, n23155, n23156, n23157, n23158, n23159,
         n23160, n23161, n23162, n23163, n23164, n23165, n23166, n23167,
         n23168, n23169, n23170, n23171, n23172, n23173, n23174, n23175,
         n23176, n23177, n23178, n23179, n23180, n23181, n23182, n23183,
         n23184, n23185, n23186, n23187, n23188, n23189, n23190, n23191,
         n23192, n23193, n23194, n23195, n23196, n23197, n23198, n23199,
         n23200, n23201, n23202, n23203, n23204, n23205, n23206, n23207,
         n23208, n23209, n23210, n23211, n23212, n23213, n23214, n23215,
         n23216, n23217, n23218, n23219, n23220, n23221, n23222, n23223,
         n23224, n23225, n23226, n23227, n23228, n23229, n23230, n23231,
         n23232, n23233, n23234, n23235, n23236, n23237, n23238, n23239,
         n23240, n23241, n23242, n23243, n23244, n23245, n23246, n23247,
         n23248, n23249, n23250, n23251, n23252, n23253, n23254, n23255,
         n23256, n23257, n23258, n23259, n23260, n23261, n23262, n23263,
         n23264, n23265, n23266, n23267, n23268, n23269, n23270, n23271,
         n23272, n23273, n23274, n23275, n23276, n23277, n23278, n23279,
         n23280, n23281, n23282, n23283, n23284, n23285, n23286, n23287,
         n23288, n23289, n23290, n23291, n23292, n23293, n23294, n23295,
         n23296, n23297, n23298, n23299, n23300, n23301, n23302, n23303,
         n23304, n23305, n23306, n23307, n23308, n23309, n23310, n23311,
         n23312, n23313, n23314, n23315, n23316, n23317, n23318, n23319,
         n23320, n23321, n23322, n23323, n23324, n23325, n23326, n23327,
         n23328, n23329, n23330, n23331, n23332, n23333, n23334, n23335,
         n23336, n23337, n23338, n23339, n23340, n23341, n23342, n23343,
         n23344, n23345, n23346, n23347, n23348, n23349, n23350, n23351,
         n23352, n23353, n23354, n23355, n23356, n23357, n23358, n23359,
         n23360, n23361, n23362, n23363, n23364, n23365, n23366, n23367,
         n23368, n23369, n23370, n23371, n23372, n23373, n23374, n23375,
         n23376, n23377, n23378, n23379, n23380, n23381, n23382, n23383,
         n23384, n23385, n23386, n23387, n23388, n23389, n23390, n23391,
         n23392, n23393, n23394, n23395, n23396, n23397, n23398, n23399,
         n23400, n23401, n23402, n23403, n23404, n23405, n23406, n23407,
         n23408, n23409, n23410, n23411, n23412, n23413, n23414, n23415,
         n23416, n23417, n23418, n23419, n23420, n23421, n23422, n23423,
         n23424, n23425, n23426, n23427, n23428, n23429, n23430, n23431,
         n23432, n23433, n23434, n23435, n23436, n23437, n23438, n23439,
         n23440, n23441, n23442, n23443, n23444, n23445, n23446, n23447,
         n23448, n23449, n23450, n23451, n23452, n23453, n23454, n23455,
         n23456, n23457, n23458, n23459, n23460, n23461, n23462, n23463,
         n23464, n23465, n23466, n23467, n23468, n23469, n23470, n23471,
         n23472, n23473, n23474, n23475, n23476, n23477, n23478, n23479,
         n23480, n23481, n23482, n23483, n23484, n23485, n23486, n23487,
         n23488, n23489, n23490, n23491, n23492, n23493, n23494, n23495,
         n23496, n23497, n23498, n23499, n23500, n23501, n23502, n23503,
         n23504, n23505, n23506, n23507, n23508, n23509, n23510, n23511,
         n23512, n23513, n23514, n23515, n23516, n23517, n23518, n23519,
         n23520, n23521, n23522, n23523, n23524, n23525, n23526, n23527,
         n23528, n23529, n23530, n23531, n23532, n23533, n23534, n23535,
         n23536, n23537, n23538, n23539, n23540, n23541, n23542, n23543,
         n23544, n23545, n23546, n23547, n23548, n23549, n23550, n23551,
         n23552, n23553, n23554, n23555, n23556, n23557, n23558, n23559,
         n23560, n23561, n23562, n23563, n23564, n23565, n23566, n23567,
         n23568, n23569, n23570, n23571, n23572, n23573, n23574, n23575,
         n23576, n23577, n23578, n23579, n23580, n23581, n23582, n23583,
         n23584, n23585, n23586, n23587, n23588, n23589, n23590, n23591,
         n23592, n23593, n23594, n23595, n23596, n23597, n23598, n23599,
         n23600, n23601, n23602, n23603, n23604, n23605, n23606, n23607,
         n23608, n23609, n23610, n23611, n23612, n23613, n23614, n23615,
         n23616, n23617, n23618, n23619, n23620, n23621, n23622, n23623,
         n23624, n23625, n23626, n23627, n23628, n23629, n23630, n23631,
         n23632, n23633, n23634, n23635, n23636, n23637, n23638, n23639,
         n23640, n23641, n23642, n23643, n23644, n23645, n23646, n23647,
         n23648, n23649, n23650, n23651, n23652, n23653, n23654, n23655,
         n23656, n23657, n23658, n23659, n23660, n23661, n23662, n23663,
         n23664, n23665, n23666, n23667, n23668, n23669, n23670, n23671,
         n23672, n23673, n23674, n23675, n23676, n23677, n23678, n23679,
         n23680, n23681, n23682, n23683, n23684, n23685, n23686, n23687,
         n23688, n23689, n23690, n23691, n23692, n23693, n23694, n23695,
         n23696, n23697, n23698, n23699, n23700, n23701, n23702, n23703,
         n23704, n23705, n23706, n23707, n23708, n23709, n23710, n23711,
         n23712, n23713, n23714, n23715, n23716, n23717, n23718, n23719,
         n23720, n23721, n23722, n23723, n23724, n23725, n23726, n23727,
         n23728, n23729, n23730, n23731, n23732, n23733, n23734, n23735,
         n23736, n23737, n23738, n23739, n23740, n23741, n23742, n23743,
         n23744, n23745, n23746, n23747, n23748, n23749, n23750, n23751,
         n23752, n23753, n23754, n23755, n23756, n23757, n23758, n23759,
         n23760, n23761, n23762, n23763, n23764, n23765, n23766, n23767,
         n23768, n23769, n23770, n23771, n23772, n23773, n23774, n23775,
         n23776, n23777, n23778, n23779, n23780, n23781, n23782, n23783,
         n23784, n23785, n23786, n23787, n23788, n23789, n23790, n23791,
         n23792, n23793, n23794, n23795, n23796, n23797, n23798, n23799,
         n23800, n23801, n23802, n23803, n23804, n23805, n23806, n23807,
         n23808, n23809, n23810, n23811, n23812, n23813, n23814, n23815,
         n23816, n23817, n23818, n23819, n23820, n23821, n23822, n23823,
         n23824, n23825, n23826, n23827, n23828, n23829, n23830, n23831,
         n23832, n23833, n23834, n23835, n23836, n23837, n23838, n23839,
         n23840, n23841, n23842, n23843, n23844, n23845, n23846, n23847,
         n23848, n23849, n23850, n23851, n23852, n23853, n23854, n23855,
         n23856, n23857, n23858, n23859, n23860, n23861, n23862, n23863,
         n23864, n23865, n23866, n23867, n23868, n23869, n23870, n23871,
         n23872, n23873, n23874, n23875, n23876, n23877, n23878, n23879,
         n23880, n23881, n23882, n23883, n23884, n23885, n23886, n23887,
         n23888, n23889, n23890, n23891, n23892, n23893, n23894, n23895,
         n23896, n23897, n23898, n23899, n23900, n23901, n23902, n23903,
         n23904, n23905, n23906, n23907, n23908, n23909, n23910, n23911,
         n23912, n23913, n23914, n23915, n23916, n23917, n23918, n23919,
         n23920, n23921, n23922, n23923, n23924, n23925, n23926, n23927,
         n23928, n23929, n23930, n23931, n23932, n23933, n23934, n23935,
         n23936, n23937, n23938, n23939, n23940, n23941, n23942, n23943,
         n23944, n23945, n23946, n23947, n23948, n23949, n23950, n23951,
         n23952, n23953, n23954, n23955, n23956, n23957, n23958, n23959,
         n23960, n23961, n23962, n23963, n23964, n23965, n23966, n23967,
         n23968, n23969, n23970, n23971, n23972, n23973, n23974, n23975,
         n23976, n23977, n23978, n23979, n23980, n23981, n23982, n23983,
         n23984, n23985, n23986, n23987, n23988, n23989, n23990, n23991,
         n23992, n23993, n23994, n23995, n23996, n23997, n23998, n23999,
         n24000, n24001, n24002, n24003, n24004, n24005, n24006, n24007,
         n24008, n24009, n24010, n24011, n24012, n24013, n24014, n24015,
         n24016, n24017, n24018, n24019, n24020, n24021, n24022, n24023,
         n24024, n24025, n24026, n24027, n24028, n24029, n24030, n24031,
         n24032, n24033, n24034, n24035, n24036, n24037, n24038, n24039,
         n24040, n24041, n24042, n24043, n24044, n24045, n24046, n24047,
         n24048, n24049, n24050, n24051, n24052, n24053, n24054, n24055,
         n24056, n24057, n24058, n24059, n24060, n24061, n24062, n24063,
         n24064, n24065, n24066, n24067, n24068, n24069, n24070, n24071,
         n24072, n24073, n24074, n24075, n24076, n24077, n24078, n24079,
         n24080, n24081, n24082, n24083, n24084, n24085, n24086, n24087,
         n24088, n24089, n24090, n24091, n24092, n24093, n24094, n24095,
         n24096, n24097, n24098, n24099, n24100, n24101, n24102, n24103,
         n24104, n24105, n24106, n24107, n24108, n24109, n24110, n24111,
         n24112, n24113, n24114, n24115, n24116, n24117, n24118, n24119,
         n24120, n24121, n24122, n24123, n24124, n24125, n24126, n24127,
         n24128, n24129, n24130, n24131, n24132, n24133, n24134, n24135,
         n24136, n24137, n24138, n24139, n24140, n24141, n24142, n24143,
         n24144, n24145, n24146, n24147, n24148, n24149, n24150, n24151,
         n24152, n24153, n24154, n24155, n24156, n24157, n24158, n24159,
         n24160, n24161, n24162, n24163, n24164, n24165, n24166, n24167,
         n24168, n24169, n24170, n24171, n24172, n24173, n24174, n24175,
         n24176, n24177, n24178, n24179, n24180, n24181, n24182, n24183,
         n24184, n24185, n24186, n24187, n24188, n24189, n24190, n24191,
         n24192, n24193, n24194, n24195, n24196, n24197, n24198, n24199,
         n24200, n24201, n24202, n24203, n24204, n24205, n24206, n24207,
         n24208, n24209, n24210, n24211, n24212, n24213, n24214, n24215,
         n24216, n24217, n24218, n24219, n24220, n24221, n24222, n24223,
         n24224, n24225, n24226, n24227, n24228, n24229, n24230, n24231,
         n24232, n24233, n24234, n24235, n24236, n24237, n24238, n24239,
         n24240, n24241, n24242, n24243, n24244, n24245, n24246, n24247,
         n24248, n24249, n24250, n24251, n24252, n24253, n24254, n24255,
         n24256, n24257, n24258, n24259, n24260, n24261, n24262, n24263,
         n24264, n24265, n24266, n24267, n24268, n24269, n24270, n24271,
         n24272, n24273, n24274, n24275, n24276, n24277, n24278, n24279,
         n24280, n24281, n24282, n24283, n24284, n24285, n24286, n24287,
         n24288, n24289, n24290, n24291, n24292, n24293, n24294, n24295,
         n24296, n24297, n24298, n24299, n24300, n24301, n24302, n24303,
         n24304, n24305, n24306, n24307, n24308, n24309, n24310, n24311,
         n24312, n24313, n24314, n24315, n24316, n24317, n24318, n24319,
         n24320, n24321, n24322, n24323, n24324, n24325, n24326, n24327,
         n24328, n24329, n24330, n24331, n24332, n24333, n24334, n24335,
         n24336, n24337, n24338, n24339, n24340, n24341, n24342, n24343,
         n24344, n24345, n24346, n24347, n24348, n24349, n24350, n24351,
         n24352, n24353, n24354, n24355, n24356, n24357, n24358, n24359,
         n24360, n24361, n24362, n24363, n24364, n24365, n24366, n24367,
         n24368, n24369, n24370, n24371, n24372, n24373, n24374, n24375,
         n24376, n24377, n24378, n24379, n24380, n24381, n24382, n24383,
         n24384, n24385, n24386, n24387, n24388, n24389, n24390, n24391,
         n24392, n24393, n24394, n24395, n24396, n24397, n24398, n24399,
         n24400, n24401, n24402, n24403, n24404, n24405, n24406, n24407,
         n24408, n24409, n24410, n24411, n24412, n24413, n24414, n24415,
         n24416, n24417, n24418, n24419, n24420, n24421, n24422, n24423,
         n24424, n24425, n24426, n24427, n24428, n24429, n24430, n24431,
         n24432, n24433, n24434, n24435, n24436, n24437, n24438, n24439,
         n24440, n24441, n24442, n24443, n24444, n24445, n24446, n24447,
         n24448, n24449, n24450, n24451, n24452, n24453, n24454, n24455,
         n24456, n24457, n24458, n24459, n24460, n24461, n24462, n24463,
         n24464, n24465, n24466, n24467, n24468, n24469, n24470, n24471,
         n24472, n24473, n24474, n24475, n24476, n24477, n24478, n24479,
         n24480, n24481, n24482, n24483, n24484, n24485, n24486, n24487,
         n24488, n24489, n24490, n24491, n24492, n24493, n24494, n24495,
         n24496, n24497, n24498, n24499, n24500, n24501, n24502, n24503,
         n24504, n24505, n24506, n24507, n24508, n24509, n24510, n24511,
         n24512, n24513, n24514, n24515, n24516, n24517, n24518, n24519,
         n24520, n24521, n24522, n24523, n24524, n24525, n24526, n24527,
         n24528, n24529, n24530, n24531, n24532, n24533, n24534, n24535,
         n24536, n24537, n24538, n24539, n24540, n24541, n24542, n24543,
         n24544, n24545, n24546, n24547, n24548, n24549, n24550, n24551,
         n24552, n24553, n24554, n24555, n24556, n24557, n24558, n24559,
         n24560, n24561, n24562, n24563, n24564, n24565, n24566, n24567,
         n24568, n24569, n24570, n24571, n24572, n24573, n24574, n24575,
         n24576, n24577, n24578, n24579, n24580, n24581, n24582, n24583,
         n24584, n24585, n24586, n24587, n24588, n24589, n24590, n24591,
         n24592, n24593, n24594, n24595, n24596, n24597, n24598, n24599,
         n24600, n24601, n24602, n24603, n24604, n24605, n24606, n24607,
         n24608, n24609, n24610, n24611, n24612, n24613, n24614, n24615,
         n24616, n24617, n24618, n24619, n24620, n24621, n24622, n24623,
         n24624, n24625, n24626, n24627, n24628, n24629, n24630, n24631,
         n24632, n24633, n24634, n24635, n24636, n24637, n24638, n24639,
         n24640, n24641, n24642, n24643, n24644, n24645, n24646, n24647,
         n24648, n24649, n24650, n24651, n24652, n24653, n24654, n24655,
         n24656, n24657, n24658, n24659, n24660, n24661, n24662, n24663,
         n24664, n24665, n24666, n24667, n24668, n24669, n24670, n24671,
         n24672, n24673, n24674, n24675, n24676, n24677, n24678, n24679,
         n24680, n24681, n24682, n24683, n24684, n24685, n24686, n24687,
         n24688, n24689, n24690, n24691, n24692, n24693, n24694, n24695,
         n24696, n24697, n24698, n24699, n24700, n24701, n24702, n24703,
         n24704, n24705, n24706, n24707, n24708, n24709, n24710, n24711,
         n24712, n24713, n24714, n24715, n24716, n24717, n24718, n24719,
         n24720, n24721, n24722, n24723, n24724, n24725, n24726, n24727,
         n24728, n24729, n24730, n24731, n24732, n24733, n24734, n24735,
         n24736, n24737, n24738, n24739, n24740, n24741, n24742, n24743,
         n24744, n24745, n24746, n24747, n24748, n24749, n24750, n24751,
         n24752, n24753, n24754, n24755, n24756, n24757, n24758, n24759,
         n24760, n24761, n24762, n24763, n24764, n24765, n24766, n24767,
         n24768, n24769, n24770, n24771, n24772, n24773, n24774, n24775,
         n24776, n24777, n24778, n24779, n24780, n24781, n24782, n24783,
         n24784, n24785, n24786, n24787, n24788, n24789, n24790, n24791,
         n24792, n24793, n24794, n24795, n24796, n24797, n24798, n24799,
         n24800, n24801, n24802, n24803, n24804, n24805, n24806, n24807,
         n24808, n24809, n24810, n24811, n24812, n24813, n24814, n24815,
         n24816, n24817, n24818, n24819, n24820, n24821, n24822, n24823,
         n24824, n24825, n24826, n24827, n24828, n24829, n24830, n24831,
         n24832, n24833, n24834, n24835, n24836, n24837, n24838, n24839,
         n24840, n24841, n24842, n24843, n24844, n24845, n24846, n24847,
         n24848, n24849, n24850, n24851, n24852, n24853, n24854, n24855,
         n24856, n24857, n24858, n24859, n24860, n24861, n24862, n24863,
         n24864, n24865, n24866, n24867, n24868, n24869, n24870, n24871,
         n24872, n24873, n24874, n24875, n24876, n24877, n24878, n24879,
         n24880, n24881, n24882, n24883, n24884, n24885, n24886, n24887,
         n24888, n24889, n24890, n24891, n24892, n24893, n24894, n24895,
         n24896, n24897, n24898, n24899, n24900, n24901, n24902, n24903,
         n24904, n24905, n24906, n24907, n24908, n24909, n24910, n24911,
         n24912, n24913, n24914, n24915, n24916, n24917, n24918, n24919,
         n24920, n24921, n24922, n24923, n24924, n24925, n24926, n24927,
         n24928, n24929, n24930, n24931, n24932, n24933, n24934, n24935,
         n24936, n24937, n24938, n24939, n24940, n24941, n24942, n24943,
         n24944, n24945, n24946, n24947, n24948, n24949, n24950, n24951,
         n24952, n24953, n24954, n24955, n24956, n24957, n24958, n24959,
         n24960, n24961, n24962, n24963, n24964, n24965, n24966, n24967,
         n24968, n24969, n24970, n24971, n24972, n24973, n24974, n24975,
         n24976, n24977, n24978, n24979, n24980, n24981, n24982, n24983,
         n24984, n24985, n24986, n24987, n24988, n24989, n24990, n24991,
         n24992, n24993, n24994, n24995, n24996, n24997, n24998, n24999,
         n25000, n25001, n25002, n25003, n25004, n25005, n25006, n25007,
         n25008, n25009, n25010, n25011, n25012, n25013, n25014, n25015,
         n25016, n25017, n25018, n25019, n25020, n25021, n25022, n25023,
         n25024, n25025, n25026, n25027, n25028, n25029, n25030, n25031,
         n25032, n25033, n25034, n25035, n25036, n25037, n25038, n25039,
         n25040, n25041, n25042, n25043, n25044, n25045, n25046, n25047,
         n25048, n25049, n25050, n25051, n25052, n25053, n25054, n25055,
         n25056, n25057, n25058, n25059, n25060, n25061, n25062, n25063,
         n25064, n25065, n25066, n25067, n25068, n25069, n25070, n25071,
         n25072, n25073, n25074, n25075, n25076, n25077, n25078, n25079,
         n25080, n25081, n25082, n25083, n25084, n25085, n25086, n25087,
         n25088, n25089, n25090, n25091, n25092, n25093, n25094, n25095,
         n25096, n25097, n25098, n25099, n25100, n25101, n25102, n25103,
         n25104, n25105, n25106, n25107, n25108, n25109, n25110, n25111,
         n25112, n25113, n25114, n25115, n25116, n25117, n25118, n25119,
         n25120, n25121, n25122, n25123, n25124, n25125, n25126, n25127,
         n25128, n25129, n25130, n25131, n25132, n25133, n25134, n25135,
         n25136, n25137, n25138, n25139, n25140, n25141, n25142, n25143,
         n25144, n25145, n25146, n25147, n25148, n25149, n25150, n25151,
         n25152, n25153, n25154, n25155, n25156, n25157, n25158, n25159,
         n25160, n25161, n25162, n25163, n25164, n25165, n25166, n25167,
         n25168, n25169, n25170, n25171, n25172, n25173, n25174, n25175,
         n25176, n25177, n25178, n25179, n25180, n25181, n25182, n25183,
         n25184, n25185, n25186, n25187, n25188, n25189, n25190, n25191,
         n25192, n25193, n25194, n25195, n25196, n25197, n25198, n25199,
         n25200, n25201, n25202, n25203, n25204, n25205, n25206, n25207,
         n25208, n25209, n25210, n25211, n25212, n25213, n25214, n25215,
         n25216, n25217, n25218, n25219, n25220, n25221, n25222, n25223,
         n25224, n25225, n25226, n25227, n25228, n25229, n25230, n25231,
         n25232, n25233, n25234, n25235, n25236, n25237, n25238, n25239,
         n25240, n25241, n25242, n25243, n25244, n25245, n25246, n25247,
         n25248, n25249, n25250, n25251, n25252, n25253, n25254, n25255,
         n25256, n25257, n25258, n25259, n25260, n25261, n25262, n25263,
         n25264, n25265, n25266, n25267, n25268, n25269, n25270, n25271,
         n25272, n25273, n25274, n25275, n25276, n25277, n25278, n25279,
         n25280, n25281, n25282, n25283, n25284, n25285, n25286, n25287,
         n25288, n25289, n25290, n25291, n25292, n25293, n25294, n25295,
         n25296, n25297, n25298, n25299, n25300, n25301, n25302, n25303,
         n25304, n25305, n25306, n25307, n25308, n25309, n25310, n25311,
         n25312, n25313, n25314, n25315, n25316, n25317, n25318, n25319,
         n25320, n25321, n25322, n25323, n25324, n25325, n25326, n25327,
         n25328, n25329, n25330, n25331, n25332, n25333, n25334, n25335,
         n25336, n25337, n25338, n25339, n25340, n25341, n25342, n25343,
         n25344, n25345, n25346, n25347, n25348, n25349, n25350, n25351,
         n25352, n25353, n25354, n25355, n25356, n25357, n25358, n25359,
         n25360, n25361, n25362, n25363, n25364, n25365, n25366, n25367,
         n25368, n25369, n25370, n25371, n25372, n25373, n25374, n25375,
         n25376, n25377, n25378, n25379, n25380, n25381, n25382, n25383,
         n25384, n25385, n25386, n25387, n25388, n25389, n25390, n25391,
         n25392, n25393, n25394, n25395, n25396, n25397, n25398, n25399,
         n25400, n25401, n25402, n25403, n25404, n25405, n25406, n25407,
         n25408, n25409, n25410, n25411, n25412, n25413, n25414, n25415,
         n25416, n25417, n25418, n25419, n25420, n25421, n25422, n25423,
         n25424, n25425, n25426, n25427, n25428, n25429, n25430, n25431,
         n25432, n25433, n25434, n25435, n25436, n25437, n25438, n25439,
         n25440, n25441, n25442, n25443, n25444, n25445, n25446, n25447,
         n25448, n25449, n25450, n25451, n25452, n25453, n25454, n25455,
         n25456, n25457, n25458, n25459, n25460, n25461, n25462, n25463,
         n25464, n25465, n25466, n25467, n25468, n25469, n25470, n25471,
         n25472, n25473, n25474, n25475, n25476, n25477, n25478, n25479,
         n25480, n25481, n25482, n25483, n25484, n25485, n25486, n25487,
         n25488, n25489, n25490, n25491, n25492, n25493, n25494, n25495,
         n25496, n25497, n25498, n25499, n25500, n25501, n25502, n25503,
         n25504, n25505, n25506, n25507, n25508, n25509, n25510, n25511,
         n25512, n25513, n25514, n25515, n25516, n25517, n25518, n25519,
         n25520, n25521, n25522, n25523, n25524, n25525, n25526, n25527,
         n25528, n25529, n25530, n25531, n25532, n25533, n25534, n25535,
         n25536, n25537, n25538, n25539, n25540, n25541, n25542, n25543,
         n25544, n25545, n25546, n25547, n25548, n25549, n25550, n25551,
         n25552, n25553, n25554, n25555, n25556, n25557, n25558, n25559,
         n25560, n25561, n25562, n25563, n25564, n25565, n25566, n25567,
         n25568, n25569, n25570, n25571, n25572, n25573, n25574, n25575,
         n25576, n25577, n25578, n25579, n25580, n25581, n25582, n25583,
         n25584, n25585, n25586, n25587, n25588, n25589, n25590, n25591,
         n25592, n25593, n25594, n25595, n25596, n25597, n25598, n25599,
         n25600, n25601, n25602, n25603, n25604, n25605, n25606, n25607,
         n25608, n25609, n25610, n25611, n25612, n25613, n25614, n25615,
         n25616, n25617, n25618, n25619, n25620, n25621, n25622, n25623,
         n25624, n25625, n25626, n25627, n25628, n25629, n25630, n25631,
         n25632, n25633, n25634, n25635, n25636, n25637, n25638, n25639,
         n25640, n25641, n25642, n25643, n25644, n25645, n25646, n25647,
         n25648, n25649, n25650, n25651, n25652, n25653, n25654, n25655,
         n25656, n25657, n25658, n25659, n25660, n25661, n25662, n25663,
         n25664, n25665, n25666, n25667, n25668, n25669, n25670, n25671,
         n25672, n25673, n25674, n25675, n25676, n25677, n25678, n25679,
         n25680, n25681, n25682, n25683, n25684, n25685, n25686, n25687,
         n25688, n25689, n25690, n25691, n25692, n25693, n25694, n25695,
         n25696, n25697, n25698, n25699, n25700, n25701, n25702, n25703,
         n25704, n25705, n25706, n25707, n25708, n25709, n25710, n25711,
         n25712, n25713, n25714, n25715, n25716, n25717, n25718, n25719,
         n25720, n25721, n25722, n25723, n25724, n25725, n25726, n25727,
         n25728, n25729, n25730, n25731, n25732, n25733, n25734, n25735,
         n25736, n25737, n25738, n25739, n25740, n25741, n25742, n25743,
         n25744, n25745, n25746, n25747, n25748, n25749, n25750, n25751,
         n25752, n25753, n25754, n25755, n25756, n25757, n25758, n25759,
         n25760, n25761, n25762, n25763, n25764, n25765, n25766, n25767,
         n25768, n25769, n25770, n25771, n25772, n25773, n25774, n25775,
         n25776, n257770, n257780, n25779, n25780, n25781, n25782, n25783,
         n25784, n25785, n25786, n25787, n25788, n25789, n25790, n25791,
         n25792, n25793, n25794, n25795, n25796, n25797, n25798, n25799,
         n25800, n25801, n25802, n25803, n25804, n25805, n25806, n25807,
         n25808, n25809, n25810, n25811, n25812, n25813, n25814, n25815,
         n25816, n25817, n25818, n25819, n25820, n25821, n25822, n25823,
         n25824, n25825, n25826, n25827, n25828, n25829, n25830, n25831,
         n25832, n25833, n25834, n25835, n25836, n25837, n25838, n25839,
         n25840, n25841, n25842, n25843, n25844, n25845, n25846, n25847,
         n25848, n25849, n25850, n25851, n25852, n25853, n25854, n25855,
         n25856, n25857, n25858, n25859, n25860, n25861, n25862, n25863,
         n25864, n25865, n25866, n25867, n25868, n25869, n25870, n25871,
         n25872, n25873, n25874, n25875, n25876, n25877, n25878, n25879,
         n25880, n25881, n25882, n25883, n25884, n25885, n25886, n25887,
         n25888, n25889, n25890, n25891, n25892, n25893, n258940, n25895,
         n25896, n25897, n25898, n25899, n25900, n25901, n25902, n25903,
         n25904, n25905, n25906, n25907, n25908, n25909, n25910, n25911,
         n25912, n25913, n25914, n25915, n25916, n25917, n25918, n25919,
         n25920, n25921, n25922, n25923, n25924, n25925, n25926, n25927,
         n25928, n25929, n25930, n25931, n25932, n25933, n25934, n25935,
         n25936, n25937, n25938, n25939, n25940, n25941, n25942, n25943,
         n25944, n25945, n25946, n25947, n25948, n25949, n25950, n25951,
         n25952, n25953, n25954, n25955, n25956, n25957, n25958, n25959,
         n25960, n25961, n25962, n25963, n25964, n25965, n25966, n25967,
         n25968, n25969, n25970, n25971, n25972, n25973, n25974, n25975,
         n25976, n25977, n25978, n25979, n25980, n25981, n25982, n25983,
         n25984, n25985, n25986, n25987, n25988, n25989, n25990, n25991,
         n25992, n25993, n25994, n25995, n25996, n25997, n25998, n25999,
         n26000, n26001, n26002, n26003, n26004, n26005, n26006, n26007,
         n26008, n26009, n26010, n26011, n26012, n26013, n26014, n26015,
         n26016, n26017, n26018, n26019, n26020, n26021, n26022, n26023,
         n26024, n26025, n26026, n26027, n26028, n26029, n26030, n26031,
         n26032, n26033, n26034, n26035, n26036, n26037, n26038, n26039,
         n26040, n26041, n26042, n26043, n26044, n26045, n26046, n26047,
         n26048, n26049, n26050, n26051, n26052, n26053, n26054, n26055,
         n26056, n26057, n26058, n26059, n26060, n26061, n26062, n26063,
         n26064, n26065, n26066, n26067, n26068, n26069, n26070, n26071,
         n26072, n26073, n26074, n26075, n26076, n26077, n26078, n26079,
         n26080, n26081, n26082, n26083, n26084, n26085, n26086, n26087,
         n26088, n26089, n26090, n26091, n26092, n26093, n26094, n26095,
         n26096, n26097, n26098, n26099, n26100, n26101, n26102, n26103,
         n26104, n26105, n26106, n26107, n26108, n26109, n26110, n26111,
         n26112, n26113, n26114, n26115, n26116, n26117, n26118, n26119,
         n26120, n26121, n26122, n26123, n26124, n26125, n26126, n26127,
         n26128, n26129, n26130, n26131, n26132, n26133, n26134, n26135,
         n26136, n26137, n26138, n26139, n26140, n26141, n26142, n26143,
         n26144, n26145, n26146, n26147, n26148, n26149, n26150, n26151,
         n26152, n26153, n26154, n26155, n26156, n26157, n26158, n26159,
         n26160, n26161, n26162, n26163, n26164, n26165, n26166, n26167,
         n26168, n26169, n26170, n26171, n26172, n26173, n26174, n26175,
         n26176, n26177, n26178, n26179, n26180, n26181, n26182, n26183,
         n26184, n26185, n26186, n26187, n26188, n26189, n26190, n26191,
         n26192, n26193, n26194, n26195, n26196, n26197, n26198, n26199,
         n26200, n26201, n26202, n26203, n26204, n26205, n26206, n26207,
         n26208, n26209, n26210, n26211, n26212, n26213, n26214, n26215,
         n26216, n26217, n26218, n26219, n26220, n26221, n26222, n26223,
         n26224, n26225, n26226, n26227, n26228, n26229, n26230, n26231,
         n26232, n26233, n26234, n26235, n26236, n26237, n26238, n26239,
         n26240, n26241, n26242, n26243, n26244, n26245, n26246, n26247,
         n26248, n26249, n26250, n26251, n26252, n26253, n26254, n26255,
         n26256, n26257, n26258, n26259, n26260, n26261, n26262, n26263,
         n26264, n26265, n26266, n26267, n26268, n26269, n26270, n26271,
         n26272, n26273, n26274, n26275, n26276, n26277, n26278, n26279,
         n26280, n26281, n26282, n26283, n26284, n26285, n26286, n26287,
         n26288, n26289, n26290, n26291, n26292, n26293, n26294, n26295,
         n26296, n26297, n26298, n26299, n26300, n26301, n26302, n26303,
         n26304, n26305, n26306, n26307, n26308, n26309, n26310, n26311,
         n26312, n26313, n26314, n26315, n26316, n26317, n26318, n26319,
         n26320, n26321, n26322, n26323, n26324, n26325, n26326, n26327,
         n26328, n26329, n26330, n26331, n26332, n26333, n26334, n26335,
         n26336, n26337, n26338, n26339, n26340, n26341, n26342, n26343,
         n26344, n26345, n26346, n26347, n26348, n26349, n26350, n26351,
         n26352, n26353, n26354, n26355, n26356, n26357, n26358, n26359,
         n26360, n26361, n26362, n26363, n26364, n26365, n26366, n26367,
         n26368, n26369, n26370, n26371, n26372, n26373, n26374, n26375,
         n26376, n26377, n26378, n26379, n26380, n26381, n26382, n26383,
         n26384, n26385, n26386, n26387, n26388, n26389, n26390, n26391,
         n26392, n26393, n26394, n26395, n26396, n26397, n26398, n26399,
         n26400, n26401, n26402, n26403, n26404, n26405, n26406, n26407,
         n26408, n26409, n26410, n26411, n26412, n26413, n26414, n26415,
         n26416, n26417, n26418, n26419, n26420, n26421, n26422, n26423,
         n26424, n26425, n26426, n26427, n26428, n26429, n26430, n26431,
         n26432, n26433, n26434, n26435, n26436, n26437, n26438, n26439,
         n26440, n26441, n26442, n26443, n26444, n26445, n26446, n26447,
         n26448, n26449, n26450, n26451, n26452, n26453, n26454, n26455,
         n26456, n26457, n26458, n26459, n26460, n26461, n26462, n26463,
         n26464, n26465, n26466, n26467, n26468, n26469, n26470, n26471,
         n26472, n26473, n26474, n26475, n26476, n26477, n26478, n26479,
         n26480, n26481, n26482, n26483, n26484, n26485, n26486, n26487,
         n26488, n26489, n26490, n26491, n26492, n26493, n26494, n26495,
         n26496, n26497, n26498, n26499, n26500, n26501, n26502, n26503,
         n26504, n26505, n26506, n26507, n26508, n26509, n26510, n26511,
         n26512, n26513, n26514, n26515, n26516, n26517, n26518, n26519,
         n26520, n26521, n26522, n26523, n26524, n26525, n26526, n26527,
         n26528, n26529, n26530, n26531, n26532, n26533, n26534, n26535,
         n26536, n26537, n26538, n26539, n26540, n26541, n26542, n26543,
         n26544, n26545, n26546, n26547, n26548, n26549, n26550, n26551,
         n26552, n26553, n26554, n26555, n26556, n26557, n26558, n26559,
         n26560, n26561, n26562, n26563, n26564, n26565, n26566, n26567,
         n26568, n26569, n26570, n26571, n26572, n26573, n26574, n26575,
         n26576, n26577, n26578, n26579, n26580, n26581, n26582, n26583,
         n26584, n26585, n26586, n26587, n26588, n26589, n26590, n26591,
         n26592, n26593, n26594, n26595, n26596, n26597, n26598, n26599,
         n26600, n26601, n26602, n26603, n26604, n26605, n26606, n26607,
         n26608, n26609, n26610, n26611, n26612, n26613, n26614, n26615,
         n26616, n26617, n26618, n26619, n26620, n26621, n26622, n26623,
         n26624, n26625, n26626, n26627, n26628, n26629, n26630, n26631,
         n26632, n26633, n26634, n26635, n26636, n26637, n26638, n26639,
         n26640, n26641, n26642, n26643, n26644, n26645, n26646, n26647,
         n26648, n26649, n26650, n26651, n26652, n26653, n26654, n26655,
         n26656, n26657, n26658, n26659, n26660, n26661, n26662, n26663,
         n26664, n26665, n26666, n26667, n26668, n26669, n26670, n26671,
         n26672, n26673, n26674, n26675, n26676, n26677, n26678, n26679,
         n26680, n26681, n26682, n26683, n26684, n26685, n26686, n26687,
         n26688, n26689, n26690, n26691, n26692, n26693, n26694, n26695,
         n26696, n26697, n26698, n26699, n26700, n26701, n26702, n26703,
         n26704, n26705, n26706, n26707, n26708, n26709, n26710, n26711,
         n26712, n26713, n26714, n26715, n26716, n26717, n26718, n26719,
         n26720, n26721, n26722, n26723, n26724, n26725, n26726, n26727,
         n26728, n26729, n26730, n26731, n26732, n26733, n26734, n26735,
         n26736, n26737, n26738, n26739, n26740, n26741, n26742, n26743,
         n26744, n26745, n26746, n26747, n26748, n26749, n26750, n26751,
         n26752, n26753, n26754, n26755, n26756, n26757, n26758, n26759,
         n26760, n26761, n26762, n26763, n26764, n26765, n26766, n26767,
         n26768, n26769, n26770, n26771, n26772, n26773, n26774, n26775,
         n26776, n26777, n26778, n26779, n26780, n26781, n26782, n26783,
         n26784, n26785, n26786, n26787, n26788, n26789, n26790, n26791,
         n26792, n26793, n26794, n26795, n26796, n26797, n26798, n26799,
         n26800, n26801, n26802, n26803, n26804, n26805, n26806, n26807,
         n26808, n26809, n26810, n26811, n26812, n26813, n26814, n26815,
         n26816, n26817, n26818, n26819, n26820, n26821, n26822, n26823,
         n26824, n26825, n26826, n26827, n26828, n26829, n26830, n26831,
         n26832, n26833, n26834, n26835, n26836, n26837, n26838, n26839,
         n26840, n26841, n26842, n26843, n26844, n26845, n26846, n26847,
         n26848, n26849, n26850, n26851, n26852, n26853, n26854, n26855,
         n26856, n26857, n26858, n26859, n26860, n26861, n26862, n26863,
         n26864, n26865, n26866, n26867, n26868, n26869, n26870, n26871,
         n26872, n26873, n26874, n26875, n26876, n26877, n26878, n26879,
         n26880, n26881, n26882, n26883, n26884, n26885, n26886, n26887,
         n26888, n26889, n26890, n26891, n26892, n26893, n26894, n26895,
         n26896, n26897, n26898, n26899, n26900, n26901, n26902, n26903,
         n26904, n26905, n26906, n26907, n26908, n26909, n26910, n26911,
         n26912, n26913, n26914, n26915, n26916, n26917, n26918, n26919,
         n26920, n26921, n26922, n26923, n26924, n26925, n26926, n26927,
         n26928, n26929, n26930, n26931, n26932, n26933, n26934, n26935,
         n26936, n26937, n26938, n26939, n26940, n26941, n26942, n26943,
         n26944, n26945, n26946, n26947, n26948, n26949, n26950, n26951,
         n26952, n26953, n26954, n26955, n26956, n26957, n26958, n26959,
         n26960, n26961, n26962, n26963, n26964, n26965, n26966, n26967,
         n26968, n26969, n26970, n26971, n26972, n26973, n26974, n26975,
         n26976, n26977, n26978, n26979, n26980, n26981, n26982, n26983,
         n26984, n26985, n26986, n26987, n26988, n26989, n26990, n26991,
         n26992, n26993, n26994, n26995, n26996, n26997, n26998, n26999,
         n27000, n27001, n27002, n27003, n27004, n27005, n27006, n27007,
         n27008, n27009, n27010, n27011, n27012, n27013, n27014, n27015,
         n27016, n27017, n27018, n27019, n27020, n27021, n27022, n27023,
         n27024, n27025, n27026, n27027, n27028, n27029, n27030, n27031,
         n27032, n27033, n27034, n27035, n27036, n27037, n27038, n27039,
         n27040, n27041, n27042, n27043, n27044, n27045, n27046, n27047,
         n27048, n27049, n27050, n27051, n27052, n27053, n27054, n27055,
         n27056, n27057, n27058, n27059, n27060, n27061, n27062, n27063,
         n27064, n27065, n27066, n27067, n27068, n27069, n27070, n27071,
         n27072, n27073, n27074, n27075, n27076, n27077, n27078, n27079,
         n27080, n27081, n27082, n27083, n27084, n27085, n27086, n27087,
         n27088, n27089, n27090, n27091, n27092, n27093, n27094, n27095,
         n27096, n27097, n27098, n27099, n27100, n27101, n27102, n27103,
         n27104, n27105, n27106, n27107, n27108, n27109, n27110, n27111,
         n27112, n27113, n27114, n27115, n27116, n27117, n27118, n27119,
         n27120, n27121, n27122, n27123, n27124, n27125, n27126, n27127,
         n27128, n27129, n27130, n27131, n27132, n27133, n27134, n27135,
         n27136, n27137, n27138, n27139, n27140, n27141, n27142, n27143,
         n27144, n27145, n27146, n27147, n27148, n27149, n27150, n27151,
         n27152, n27153, n27154, n27155, n27156, n27157, n27158, n27159,
         n27160, n27161, n27162, n27163, n27164, n27165, n27166, n27167,
         n27168, n27169, n27170, n27171, n27172, n27173, n27174, n27175,
         n27176, n27177, n27178, n27179, n27180, n27181, n27182, n27183,
         n27184, n27185, n27186, n27187, n27188, n27189, n27190, n27191,
         n27192, n27193, n27194, n27195, n27196, n27197, n27198, n27199,
         n27200, n27201, n27202, n27203, n27204, n27205, n27206, n27207,
         n27208, n27209, n27210, n27211, n27212, n27213, n27214, n27215,
         n27216, n27217, n27218, n27219, n27220, n27221, n27222, n27223,
         n27224, n27225, n27226, n27227, n27228, n27229, n27230, n27231,
         n27232, n27233, n27234, n27235, n27236, n27237, n27238, n27239,
         n27240, n27241, n27242, n27243, n27244, n27245, n27246, n27247,
         n27248, n27249, n27250, n27251, n27252, n27253, n27254, n27255,
         n27256, n27257, n27258, n27259, n27260, n27261, n27262, n27263,
         n27264, n27265, n27266, n27267, n27268, n27269, n27270, n27271,
         n27272, n27273, n27274, n27275, n27276, n27277, n27278, n27279,
         n27280, n27281, n27282, n27283, n27284, n27285, n27286, n27287,
         n27288, n27289, n27290, n27291, n27292, n27293, n27294, n27295,
         n27296, n27297, n27298, n27299, n27300, n27301, n27302, n27303,
         n27304, n27305, n27306, n27307, n27308, n27309, n27310, n27311,
         n27312, n27313, n27314, n27315, n27316, n27317, n27318, n27319,
         n27320, n27321, n27322, n27323, n27324, n27325, n27326, n27327,
         n27328, n27329, n27330, n27331, n27332, n27333, n27334, n27335,
         n27336, n27337, n27338, n27339, n27340, n27341, n27342, n27343,
         n27344, n27345, n27346, n27347, n27348, n27349, n27350, n27351,
         n27352, n27353, n27354, n27355, n27356, n27357, n27358, n27359,
         n27360, n27361, n27362, n27363, n27364, n27365, n27366, n27367,
         n27368, n27369, n27370, n27371, n27372, n27373, n27374, n27375,
         n27376, n27377, n27378, n27379, n27380, n27381, n27382, n27383,
         n27384, n27385, n27386, n27387, n27388, n27389, n27390, n27391,
         n27392, n27393, n27394, n27395, n27396, n27397, n27398, n27399,
         n27400, n27401, n27402, n27403, n27404, n27405, n27406, n27407,
         n27408, n27409, n27410, n27411, n27412, n27413, n27414, n27415,
         n27416, n27417, n27418, n27419, n27420, n27421, n27422, n27423,
         n27424, n27425, n27426, n27427, n27428, n27429, n27430, n27431,
         n27432, n27433, n27434, n27435, n27436, n27437, n27438, n27439,
         n27440, n27441, n27442, n27443, n27444, n27445, n27446, n27447,
         n27448, n27449, n27450, n27451, n27452, n27453, n27454, n27455,
         n27456, n27457, n27458, n27459, n27460, n27461, n27462, n27463,
         n27464, n27465, n27466, n27467, n27468, n27469, n27470, n27471,
         n27472, n27473, n27474, n27475, n27476, n27477, n27478, n27479,
         n27480, n27481, n27482, n27483, n27484, n27485, n27486, n27487,
         n27488, n27489, n27490, n27491, n27492, n27493, n27494, n27495,
         n27496, n27497, n27498, n27499, n27500, n27501, n27502, n27503,
         n27504, n27505, n27506, n27507, n27508, n27509, n27510, n27511,
         n27512, n27513, n27514, n27515, n27516, n27517, n27518, n27519,
         n27520, n27521, n27522, n27523, n27524, n27525, n27526, n27527,
         n27528, n27529, n27530, n27531, n27532, n27533, n27534, n27535,
         n27536, n27537, n27538, n27539, n27540, n27541, n27542, n27543,
         n27544, n27545, n27546, n27547, n27548, n27549, n27550, n27551,
         n27552, n27553, n27554, n27555, n27556, n27557, n27558, n27559,
         n27560, n27561, n27562, n27563, n27564, n27565, n27566, n27567,
         n27568, n27569, n27570, n27571, n27572, n27573, n27574, n27575,
         n27576, n27577, n27578, n27579, n27580, n27581, n27582, n27583,
         n27584, n27585, n27586, n27587, n27588, n27589, n27590, n27591,
         n27592, n27593, n27594, n27595, n27596, n27597, n27598, n27599,
         n27600, n27601, n27602, n27603, n27604, n27605, n27606, n27607,
         n27608, n27609, n27610, n27611, n27612, n27613, n27614, n27615,
         n27616, n27617, n27618, n27619, n27620, n27621, n27622, n27623,
         n27624, n27625, n27626, n27627, n27628, n27629, n27630, n27631,
         n27632, n27633, n27634, n27635, n27636, n27637, n27638, n27639,
         n27640, n27641, n27642, n27643, n27644, n27645, n27646, n27647,
         n27648, n27649, n27650, n27651, n27652, n27653, n27654, n27655,
         n27656, n27657, n27658, n27659, n27660, n27661, n27662, n27663,
         n27664, n27665, n27666, n27667, n27668, n27669, n27670, n27671,
         n27672, n27673, n27674, n27675, n27676, n27677, n27678, n27679,
         n27680, n27681, n27682, n27683, n27684, n27685, n27686, n27687,
         n27688, n27689, n27690, n27691, n27692, n27693, n27694, n27695,
         n27696, n27697, n27698, n27699, n27700, n27701, n27702, n27703,
         n27704, n27705, n27706, n27707, n27708, n27709, n27710, n27711,
         n27712, n27713, n27714, n27715, n27716, n27717, n27718, n27719,
         n27720, n27721, n27722, n27723, n27724, n27725, n27726, n27727,
         n27728, n27729, n27730, n27731, n27732, n27733, n27734, n27735,
         n27736, n27737, n27738, n27739, n27740, n27741, n27742, n27743,
         n27744, n27745, n27746, n27747, n27748, n27749, n27750, n27751,
         n27752, n27753, n27754, n27755, n27756, n27757, n27758, n27759,
         n27760, n27761, n27762, n27763, n27764, n27765, n27766, n27767,
         n27768, n27769, n27770, n27771, n27772, n27773, n27774, n27775,
         n27776, n27777, n27778, n27779, n27780, n27781, n27782, n27783,
         n27784, n27785, n27786, n27787, n27788, n27789, n27790, n27791,
         n27792, n27793, n27794, n27795, n27796, n27797, n27798, n27799,
         n27800, n27801, n27802, n27803, n27804, n27805, n27806, n27807,
         n27808, n27809, n27810, n27811, n27812, n27813, n27814, n27815,
         n27816, n27817, n27818, n27819, n27820, n27821, n27822, n27823,
         n27824, n27825, n27826, n27827, n27828, n27829, n27830, n27831,
         n27832, n27833, n27834, n27835, n27836, n27837, n27838, n27839,
         n27840, n27841, n27842, n27843, n27844, n27845, n27846, n27847,
         n27848, n27849, n27850, n27851, n27852, n27853, n27854, n27855,
         n27856, n27857, n27858, n27859, n27860, n27861, n27862, n27863,
         n27864, n27865, n27866, n27867, n27868, n27869, n27870, n27871,
         n27872, n27873, n27874, n27875, n27876, n27877, n27878, n27879,
         n27880, n27881, n27882, n27883, n27884, n27885, n27886, n27887,
         n27888, n27889, n27890, n27891, n27892, n27893, n27894, n27895,
         n27896, n27897, n27898, n27899, n27900, n27901, n27902, n27903,
         n27904, n27905, n27906, n27907, n27908, n27909, n27910, n27911,
         n27912, n27913, n27914, n27915, n27916, n27917, n27918, n27919,
         n27920, n27921, n27922, n27923, n27924, n27925, n27926, n27927,
         n27928, n27929, n27930, n27931, n27932, n27933, n27934, n27935,
         n27936, n27937, n27938, n27939, n27940, n27941, n27942, n27943,
         n27944, n27945, n27946, n27947, n27948, n27949, n27950, n27951,
         n27952, n27953, n27954, n27955, n27956, n27957, n27958, n27959,
         n27960, n27961, n27962, n27963, n27964, n27965, n27966, n27967,
         n27968, n27969, n27970, n27971, n27972, n27973, n27974, n27975,
         n27976, n27977, n27978, n27979, n27980, n27981, n27982, n27983,
         n27984, n27985, n27986, n27987, n27988, n27989, n27990, n27991,
         n27992, n27993, n27994, n27995, n27996, n27997, n27998, n27999,
         n28000, n28001, n28002, n28003, n28004, n28005, n28006, n28007,
         n28008, n28009, n28010, n28011, n28012, n28013, n28014, n28015,
         n28016, n28017, n28018, n28019, n28020, n28021, n28022, n28023,
         n28024, n28025, n28026, n28027, n28028, n28029, n28030, n28031,
         n28032, n28033, n28034, n28035, n28036, n28037, n28038, n28039,
         n28040, n28041, n28042, n28043, n28044, n28045, n28046, n28047,
         n28048, n28049, n28050, n28051, n28052, n28053, n28054, n28055,
         n28056, n28057, n28058, n28059, n28060, n28061, n28062, n28063,
         n28064, n28065, n28066, n28067, n28068, n28069, n28070, n28071,
         n28072, n28073, n28074, n28075, n28076, n28077, n28078, n28079,
         n28080, n28081, n28082, n28083, n28084, n28085, n28086, n28087,
         n28088, n28089, n28090, n28091, n28092, n28093, n28094, n28095,
         n28096, n28097, n28098, n28099, n28100, n28101, n28102, n28103,
         n28104, n28105, n28106, n28107, n28108, n28109, n28110, n28111,
         n28112, n28113, n28114, n28115, n28116, n28117, n28118, n28119,
         n28120, n28121, n28122, n28123, n28124, n28125, n28126, n28127,
         n28128, n28129, n28130, n28131, n28132, n28133, n28134, n28135,
         n28136, n28137, n28138, n28139, n28140, n28141, n28142, n28143,
         n28144, n28145, n28146, n28147, n28148, n28149, n28150, n28151,
         n28152, n28153, n28154, n28155, n28156, n28157, n28158, n28159,
         n28160, n28161, n28162, n28163, n28164, n28165, n28166, n28167,
         n28168, n28169, n28170, n28171, n28172, n28173, n28174, n28175,
         n28176, n28177, n28178, n28179, n28180, n28181, n28182, n28183,
         n28184, n28185, n28186, n28187, n28188, n28189, n28190, n28191,
         n28192, n28193, n28194, n28195, n28196, n28197, n28198, n28199,
         n28200, n28201, n28202, n28203, n28204, n28205, n28206, n28207,
         n28208, n28209, n28210, n28211, n28212, n28213, n28214, n28215,
         n28216, n28217, n28218, n28219, n28220, n28221, n28222, n28223,
         n28224, n28225, n28226, n28227, n28228, n28229, n28230, n28231,
         n28232, n28233, n28234, n28235, n28236, n28237, n28238, n28239,
         n28240, n28241, n28242, n28243, n28244, n28245, n28246, n28247,
         n28248, n28249, n28250, n28251, n28252, n28253, n28254, n28255,
         n28256, n28257, n28258, n28259, n28260, n28261, n28262, n28263,
         n28264, n28265, n28266, n28267, n28268, n28269, n28270, n28271,
         n28272, n28273, n28274, n28275, n28276, n28277, n28278, n28279,
         n28280, n28281, n28282, n28283, n28284, n28285, n28286, n28287,
         n28288, n28289, n28290, n28291, n28292, n28293, n28294, n28295,
         n28296, n28297, n28298, n28299, n28300, n28301, n28302, n28303,
         n28304, n28305, n28306, n28307, n28308, n28309, n28310, n28311,
         n28312, n28313, n28314, n28315, n28316, n28317, n28318, n28319,
         n28320, n28321, n28322, n28323, n28324, n28325, n28326, n28327,
         n28328, n28329, n28330, n28331, n28332, n28333, n28334, n28335,
         n28336, n28337, n28338, n28339, n28340, n28341, n28342, n28343,
         n28344, n28345, n28346, n28347, n28348, n28349, n28350, n28351,
         n28352, n28353, n28354, n28355, n28356, n28357, n28358, n28359,
         n28360, n28361, n28362, n28363, n28364, n28365, n28366, n28367,
         n28368, n28369, n28370, n28371, n28372, n28373, n28374, n28375,
         n28376, n28377, n28378, n28379, n28380, n28381, n28382, n28383,
         n28384, n28385, n28386, n28387, n28388, n28389, n28390, n28391,
         n28392, n28393, n28394, n28395, n28396, n28397, n28398, n28399,
         n28400, n28401, n28402, n28403, n28404, n28405, n28406, n28407,
         n28408, n28409, n28410, n28411, n28412, n28413, n28414, n28415,
         n28416, n28417, n28418, n28419, n28420, n28421, n28422, n28423,
         n28424, n28425, n28426, n28427, n28428, n28429, n28430, n28431,
         n28432, n28433, n28434, n28435, n28436, n28437, n28438, n28439,
         n28440, n28441, n28442, n28443, n28444, n28445, n28446, n28447,
         n28448, n28449, n28450, n28451, n28452, n28453, n28454, n28455,
         n28456, n28457, n28458, n28459, n28460, n28461, n28462, n28463,
         n28464, n28465, n28466, n28467, n28468, n28469, n28470, n28471,
         n28472, n28473, n28474, n28475, n28476, n28477, n28478, n28479,
         n28480, n28481, n28482, n28483, n28484, n28485, n28486, n28487,
         n28488, n28489, n28490, n28491, n28492, n28493, n28494, n28495,
         n28496, n28497, n28498, n28499, n28500, n28501, n28502, n28503,
         n28504, n28505, n28506, n28507, n28508, n28509, n28510, n28511,
         n28512, n28513, n28514, n28515, n28516, n28517, n28518, n28519,
         n28520, n28521, n28522, n28523, n28524, n28525, n28526, n28527,
         n28528, n28529, n28530, n28531, n28532, n28533, n28534, n28535,
         n28536, n28537, n28538, n28539, n28540, n28541, n28542, n28543,
         n28544, n28545, n28546, n28547, n28548, n28549, n28550, n28551,
         n28552, n28553, n28554, n28555, n28556, n28557, n28558, n28559,
         n28560, n28561, n28562, n28563, n28564, n28565, n28566, n28567,
         n28568, n28569, n28570, n28571, n28572, n28573, n28574, n28575,
         n28576, n28577, n28578, n28579, n28580, n28581, n28582, n28583,
         n28584, n28585, n28586, n28587, n28588, n28589, n28590, n28591,
         n28592, n28593, n28594, n28595, n28596, n28597, n28598, n28599,
         n28600, n28601, n28602, n28603, n28604, n28605, n28606, n28607,
         n28608, n28609, n28610, n28611, n28612, n28613, n28614, n28615,
         n28616, n28617, n28618, n28619, n28620, n28621, n28622, n28623,
         n28624, n28625, n28626, n28627, n28628, n28629, n28630, n28631,
         n28632, n28633, n28634, n28635, n28636, n28637, n28638, n28639,
         n28640, n28641, n28642, n28643, n28644, n28645, n28646, n28647,
         n28648, n28649, n28650, n28651, n28652, n28653, n28654, n28655,
         n28656, n28657, n28658, n28659, n28660, n28661, n28662, n28663,
         n28664, n28665, n28666, n28667, n28668, n28669, n28670, n28671,
         n28672, n28673, n28674, n28675, n28676, n28677, n28678, n28679,
         n28680, n28681, n28682, n28683, n28684, n28685, n28686, n28687,
         n28688, n28689, n28690, n28691, n28692, n28693, n28694, n28695,
         n28696, n28697, n28698, n28699, n28700, n28701, n28702, n28703,
         n28704, n28705, n28706, n28707, n28708, n28709, n28710, n28711,
         n28712, n28713, n28714, n28715, n28716, n28717, n28718, n28719,
         n28720, n28721, n28722, n28723, n28724, n28725, n28726, n28727,
         n28728, n28729, n28730, n28731, n28732, n28733, n28734, n28735,
         n28736, n28737, n28738, n28739, n28740, n28741, n28742, n28743,
         n28744, n28745, n28746, n28747, n28748, n28749, n28750, n28751,
         n28752, n28753, n28754, n28755, n28756, n28757, n28758, n28759,
         n28760, n28761, n28762, n28763, n28764, n28765, n28766, n28767,
         n28768, n28769, n28770, n28771, n28772, n28773, n28774, n28775,
         n28776, n28777, n28778, n28779, n28780, n28781, n28782, n28783,
         n28784, n28785, n28786, n28787, n28788, n28789, n28790, n28791,
         n28792, n28793, n28794, n28795, n28796, n28797, n28798, n28799,
         n28800, n28801, n28802, n28803, n28804, n28805, n28806, n28807,
         n28808, n28809, n28810, n28811, n28812, n28813, n28814, n28815,
         n28816, n28817, n28818, n28819, n28820, n28821, n28822, n28823,
         n28824, n28825, n28826, n28827, n28828, n28829, n28830, n28831,
         n28832, n28833, n28834, n28835, n28836, n28837, n28838, n28839,
         n28840, n28841, n28842, n28843, n28844, n28845, n28846, n28847,
         n28848, n28849, n28850, n28851, n28852, n28853, n28854, n28855,
         n28856, n28857, n28858, n28859, n28860, n28861, n28862, n28863,
         n28864, n28865, n28866, n28867, n28868, n28869, n28870, n28871,
         n28872, n28873, n28874, n28875, n28876, n28877, n28878, n28879,
         n28880, n28881, n28882, n28883, n28884, n28885, n28886, n28887,
         n28888, n28889, n28890, n28891, n28892, n28893, n28894, n28895,
         n28896, n28897, n28898, n28899, n28900, n28901, n28902, n28903,
         n28904, n28905, n28906, n28907, n28908, n28909, n28910, n28911,
         n28912, n28913, n28914, n28915, n28916, n28917, n28918, n28919,
         n28920, n28921, n28922, n28923, n28924, n28925, n28926, n28927,
         n28928, n28929, n28930, n28931, n28932, n28933, n28934, n28935,
         n28936, n28937, n28938, n28939, n28940, n28941, n28942, n28943,
         n28944, n28945, n28946, n28947, n28948, n28949, n28950, n28951,
         n28952, n28953, n28954, n28955, n28956, n28957, n28958, n28959,
         n28960, n28961, n28962, n28963, n28964, n28965, n28966, n28967,
         n28968, n28969, n28970, n28971, n28972, n28973, n28974, n28975,
         n28976, n28977, n28978, n28979, n28980, n28981, n28982, n28983,
         n28984, n28985, n28986, n28987, n28988, n28989, n28990, n28991,
         n28992, n28993, n28994, n28995, n28996, n28997, n28998, n28999,
         n29000, n29001, n29002, n29003, n29004, n29005, n29006, n29007,
         n29008, n29009, n29010, n29011, n29012, n29013, n29014, n29015,
         n29016, n29017, n29018, n29019, n29020, n29021, n29022, n29023,
         n29024, n29025, n29026, n29027, n29028, n29029, n29030, n29031,
         n29032, n29033, n29034, n29035, n29036, n29037, n29038, n29039,
         n29040, n29041, n29042, n29043, n29044, n29045, n29046, n29047,
         n29048, n29049, n29050, n29051, n29052, n29053, n29054, n29055,
         n29056, n29057, n29058, n29059, n29060, n29061, n29062, n29063,
         n29064, n29065, n29066, n29067, n29068, n29069, n29070, n29071,
         n29072, n29073, n29074, n29075, n29076, n29077, n29078, n29079,
         n29080, n29081, n29082, n29083, n29084, n29085, n29086, n29087,
         n29088, n29089, n29090, n29091, n29092, n29093, n29094, n29095,
         n29096, n29097, n29098, n29099, n29100, n29101, n29102, n29103,
         n29104, n29105, n29106, n29107, n29108, n29109, n29110, n29111,
         n29112, n29113, n29114, n29115, n29116, n29117, n29118, n29119,
         n29120, n29121, n29122, n29123, n29124, n29125, n29126, n29127,
         n29128, n29129, n29130, n29131, n29132, n29133, n29134, n29135,
         n29136, n29137, n29138, n29139, n29140, n29141, n29142, n29143,
         n29144, n29145, n29146, n29147, n29148, n29149, n29150, n29151,
         n29152, n29153, n29154, n29155, n29156, n29157, n29158, n29159,
         n29160, n29161, n29162, n29163, n29164, n29165, n29166, n29167,
         n29168, n29169, n29170, n29171, n29172, n29173, n29174, n29175,
         n29176, n29177, n29178, n29179, n29180, n29181, n29182, n29183,
         n29184, n29185, n29186, n29187, n29188, n29189, n29190, n29191,
         n29192, n29193, n29194, n29195, n29196, n29197, n29198, n29199,
         n29200, n29201, n29202, n29203, n29204, n29205, n29206, n29207,
         n29208, n29209, n29210, n29211, n29212, n29213, n29214, n29215,
         n29216, n29217, n29218, n29219, n29220, n29221, n29222, n29223,
         n29224, n29225, n29226, n29227, n29228, n29229, n29230, n29231,
         n29232, n29233, n29234, n29235, n29236, n29237, n29238, n29239,
         n29240, n29241, n29242, n29243, n29244, n29245, n29246, n29247,
         n29248, n29249, n29250, n29251, n29252, n29253, n29254, n29255,
         n29256, n29257, n29258, n29259, n29260, n29261, n29262, n29263,
         n29264, n29265, n29266, n29267, n29268, n29269, n29270, n29271,
         n29272, n29273, n29274, n29275, n29276, n29277, n29278, n29279,
         n29280, n29281, n29282, n29283, n29284, n29285, n29286, n29287,
         n29288, n29289, n29290, n29291, n29292, n29293, n29294, n29295,
         n29296, n29297, n29298, n29299, n29300, n29301, n29302, n29303,
         n29304, n29305, n29306, n29307, n29308, n29309, n29310, n29311,
         n29312, n29313, n29314, n29315, n29316, n29317, n29318, n29319,
         n29320, n29321, n29322, n29323, n29324, n29325, n29326, n29327,
         n29328, n29329, n29330, n29331, n29332, n29333, n29334, n29335,
         n29336, n29337, n29338, n29339, n29340, n29341, n29342, n29343,
         n29344, n29345, n29346, n29347, n29348, n29349, n29350, n29351,
         n29352, n29353, n29354, n29355, n29356, n29357, n29358, n29359,
         n29360, n29361, n29362, n29363, n29364, n29365, n29366, n29367,
         n29368, n29369, n29370, n29371, n29372, n29373, n29374, n29375,
         n29376, n29377, n29378, n29379, n29380, n29381, n29382, n29383,
         n29384, n29385, n29386, n29387, n29388, n29389, n29390, n29391,
         n29392, n29393, n29394, n29395, n29396, n29397, n29398, n29399,
         n29400, n29401, n29402, n29403, n29404, n29405, n29406, n29407,
         n29408, n29409, n29410, n29411, n29412, n29413, n29414, n29415,
         n29416, n29417, n29418, n29419, n29420, n29421, n29422, n29423,
         n29424, n29425, n29426, n29427, n29428, n29429, n29430, n29431,
         n29432, n29433, n29434, n29435, n29436, n29437, n29438, n29439,
         n29440, n29441, n29442, n29443, n29444, n29445, n29446, n29447,
         n29448, n29449, n29450, n29451, n29452, n29453, n29454, n29455,
         n29456, n29457, n29458, n29459, n29460, n29461, n29462, n29463,
         n29464, n29465, n29466, n29467, n29468, n29469, n29470, n29471,
         n29472, n29473, n29474, n29475, n29476, n29477, n29478, n29479,
         n29480, n29481, n29482, n29483, n29484, n29485, n29486, n29487,
         n29488, n29489, n29490, n29491, n29492, n29493, n29494, n29495,
         n29496, n29497, n29498, n29499, n29500, n29501, n29502, n29503,
         n29504, n29505, n29506, n29507, n29508, n29509, n29510, n29511,
         n29512, n29513, n29514, n29515, n29516, n29517, n29518, n29519,
         n29520, n29521, n29522, n29523, n29524, n29525, n29526, n29527,
         n29528, n29529, n29530, n29531, n29532, n29533, n29534, n29535,
         n29536, n29537, n29538, n29539, n29540, n29541, n29542, n29543,
         n29544, n29545, n29546, n29547, n29548, n29549, n29550, n29551,
         n29552, n29553, n29554, n29555, n29556, n29557, n29558, n29559,
         n29560, n29561, n29562, n29563, n29564, n29565, n29566, n29567,
         n29568, n29569, n29570, n29571, n29572, n29573, n29574, n29575,
         n29576, n29577, n29578, n29579, n29580, n29581, n29582, n29583,
         n29584, n29585, n29586, n29587, n29588, n29589, n29590, n29591,
         n29592, n29593, n29594, n29595, n29596, n29597, n29598, n29599,
         n29600, n29601, n29602, n29603, n29604, n29605, n29606, n29607,
         n29608, n29609, n29610, n29611, n29612, n29613, n29614, n29615,
         n29616, n29617, n29618, n29619, n29620, n29621, n29622, n29623,
         n29624, n29625, n29626, n29627, n29628, n29629, n29630, n29631,
         n29632, n29633, n29634, n29635, n29636, n29637, n29638, n29639,
         n29640, n29641, n29642, n29643, n29644, n29645, n29646, n29647,
         n29648, n29649, n29650, n29651, n29652, n29653, n29654, n29655,
         n29656, n29657, n29658, n29659, n29660, n29661, n29662, n29663,
         n29664, n29665, n29666, n29667, n29668, n29669, n29670, n29671,
         n29672, n29673, n29674, n29675, n29676, n29677, n29678, n29679,
         n29680, n29681, n29682, n29683, n29684, n29685, n29686, n29687,
         n29688, n29689, n29690, n29691, n29692, n29693, n29694, n29695,
         n29696, n29697, n29698, n29699, n29700, n29701, n29702, n29703,
         n29704, n29705, n29706, n29707, n29708, n29709, n29710, n29711,
         n29712, n29713, n29714, n29715, n29716, n29717, n29718, n29719,
         n29720, n29721, n29722, n29723, n29724, n29725, n29726, n29727,
         n29728, n29729, n29730, n29731, n29732, n29733, n29734, n29735,
         n29736, n29737, n29738, n29739, n29740, n29741, n29742, n29743,
         n29744, n29745, n29746, n29747, n29748, n29749, n29750, n29751,
         n29752, n29753, n29754, n29755, n29756, n29757, n29758, n29759,
         n29760, n29761, n29762, n29763, n29764, n29765, n29766, n29767,
         n29768, n29769, n29770, n29771, n29772, n29773, n29774, n29775,
         n29776, n29777, n29778, n29779, n29780, n29781, n29782, n29783,
         n29784, n29785, n29786, n29787, n29788, n29789, n29790, n29791,
         n29792, n29793, n29794, n29795, n29796, n29797, n29798, n29799,
         n29800, n29801, n29802, n29803, n29804, n29805, n29806, n29807,
         n29808, n29809, n29810, n29811, n29812, n29813, n29814, n29815,
         n29816, n29817, n29818, n29819, n29820, n29821, n29822, n29823,
         n29824, n29825, n29826, n29827, n29828, n29829, n29830, n29831,
         n29832, n29833, n29834, n29835, n29836, n29837, n29838, n29839,
         n29840, n29841, n29842, n29843, n29844, n29845, n29846, n29847,
         n29848, n29849, n29850, n29851, n29852, n29853, n29854, n29855,
         n29856, n29857, n29858, n29859, n29860, n29861, n29862, n29863,
         n29864, n29865, n29866, n29867, n29868, n29869, n29870, n29871,
         n29872, n29873, n29874, n29875, n29876, n29877, n29878, n29879,
         n29880, n29881, n29882, n29883, n29884, n29885, n29886, n29887,
         n29888, n29889, n29890, n29891, n29892, n29893, n29894, n29895,
         n29896, n29897, n29898, n29899, n29900, n29901, n29902, n29903,
         n29904, n29905, n29906, n29907, n29908, n29909, n29910, n29911,
         n29912, n29913, n29914, n29915, n29916, n29917, n29918, n29919,
         n29920, n29921, n29922, n29923, n29924, n29925, n29926, n29927,
         n29928, n29929, n29930, n29931, n29932, n29933, n29934, n29935,
         n29936, n29937, n29938, n29939, n29940, n29941, n29942, n29943,
         n29944, n29945, n29946, n29947, n29948, n29949, n29950, n29951,
         n29952, n29953, n29954, n29955, n29956, n29957, n29958, n29959,
         n29960, n29961, n29962, n29963, n29964, n29965, n29966, n29967,
         n29968, n29969, n29970, n29971, n29972, n29973, n29974, n29975,
         n29976, n29977, n29978, n29979, n29980, n29981, n29982, n29983,
         n29984, n29985, n29986, n29987, n29988, n29989, n29990, n29991,
         n29992, n29993, n29994, n29995, n29996, n29997, n29998, n29999,
         n30000, n30001, n30002, n30003, n30004, n30005, n30006, n30007,
         n30008, n30009, n30010, n30011, n30012, n30013, n30014, n30015,
         n30016, n30017, n30018, n30019, n30020, n30021, n30022, n30023,
         n30024, n30025, n30026, n30027, n30028, n30029, n30030, n30031,
         n30032, n30033, n30034, n30035, n30036, n30037, n30038, n30039,
         n30040, n30041, n30042, n30043, n30044, n30045, n30046, n30047,
         n30048, n30049, n30050, n30051, n30052, n30053, n30054, n30055,
         n30056, n30057, n30058, n30059, n30060, n30061, n30062, n30063,
         n30064, n30065, n30066, n30067, n30068, n30069, n30070, n30071,
         n30072, n30073, n30074, n30075, n30076, n30077, n30078, n30079,
         n30080, n30081, n30082, n30083, n30084, n30085, n30086, n30087,
         n30088, n30089, n30090, n30091, n30092, n30093, n30094, n30095,
         n30096, n30097, n30098, n30099, n30100, n30101, n30102, n30103,
         n30104, n30105, n30106, n30107, n30108, n30109, n30110, n30111,
         n30112, n30113, n30114, n30115, n30116, n30117, n30118, n30119,
         n30120, n30121, n30122, n30123, n30124, n30125, n30126, n30127,
         n30128, n30129, n30130, n30131, n30132, n30133, n30134, n30135,
         n30136, n30137, n30138, n30139, n30140, n30141, n30142, n30143,
         n30144, n30145, n30146, n30147, n30148, n30149, n30150, n30151,
         n30152, n30153, n30154, n30155, n30156, n30157, n30158, n30159,
         n30160, n30161, n30162, n30163, n30164, n30165, n30166, n30167,
         n30168, n30169, n30170, n30171, n30172, n30173, n30174, n30175,
         n30176, n30177, n30178, n30179, n30180, n30181, n30182, n30183,
         n30184, n30185, n30186, n30187, n30188, n30189, n30190, n30191,
         n30192, n30193, n30194, n30195, n30196, n30197, n30198, n30199,
         n30200, n30201, n30202, n30203, n30204, n30205, n30206, n30207,
         n30208, n30209, n30210, n30211, n30212, n30213, n30214, n30215,
         n30216, n30217, n30218, n30219, n30220, n30221, n30222, n30223,
         n30224, n30225, n30226, n30227, n30228, n30229, n30230, n30231,
         n30232, n30233, n30234, n30235, n30236, n30237, n30238, n30239,
         n30240, n30241, n30242, n30243, n30244, n30245, n30246, n30247,
         n30248, n30249, n30250, n30251, n30252, n30253, n30254, n30255,
         n30256, n30257, n30258, n30259, n30260, n30261, n30262, n30263,
         n30264, n30265, n30266, n30267, n30268, n30269, n30270, n30271,
         n30272, n30273, n30274, n30275, n30276, n30277, n30278, n30279,
         n30280, n30281, n30282, n30283, n30284, n30285, n30286, n30287,
         n30288, n30289, n30290, n30291, n30292, n30293, n30294, n30295,
         n30296, n30297, n30298, n30299, n30300, n30301, n30302, n30303,
         n30304, n30305, n30306, n30307, n30308, n30309, n30310, n30311,
         n30312, n30313, n30314, n30315, n30316, n30317, n30318, n30319,
         n30320, n30321, n30322, n30323, n30324, n30325, n30326, n30327,
         n30328, n30329, n30330, n30331, n30332, n30333, n30334, n30335,
         n30336, n30337, n30338, n30339, n30340, n30341, n30342, n30343,
         n30344, n30345, n30346, n30347, n30348, n30349, n30350, n30351,
         n30352, n30353, n30354, n30355, n30356, n30357, n30358, n30359,
         n30360, n30361, n30362, n30363, n30364, n30365, n30366, n30367,
         n30368, n30369, n30370, n30371, n30372, n30373, n30374, n30375,
         n30376, n30377, n30378, n30379, n30380, n30381, n30382, n30383,
         n30384, n30385, n30386, n30387, n30388, n30389, n30390, n30391,
         n30392, n30393, n30394, n30395, n30396, n30397, n30398, n30399,
         n30400, n30401, n30402, n30403, n30404, n30405, n30406, n30407,
         n30408, n30409, n30410, n30411, n30412, n30413, n30414, n30415,
         n30416, n30417, n30418, n30419, n30420, n30421, n30422, n30423,
         n30424, n30425, n30426, n30427, n30428, n30429, n30430, n30431,
         n30432, n30433, n30434, n30435, n30436, n30437, n30438, n30439,
         n30440, n30441, n30442, n30443, n30444, n30445, n30446, n30447,
         n30448, n30449, n30450, n30451, n30452, n30453, n30454, n30455,
         n30456, n30457, n30458, n30459, n30460, n30461, n30462, n30463,
         n30464, n30465, n30466, n30467, n30468, n30469, n30470, n30471,
         n30472, n30473, n30474, n30475, n30476, n30477, n30478, n30479,
         n30480, n30481, n30482, n30483, n30484, n30485, n30486, n30487,
         n30488, n30489, n30490, n30491, n30492, n30493, n30494, n30495,
         n30496, n30497, n30498, n30499, n30500, n30501, n30502, n30503,
         n30504, n30505, n30506, n30507, n30508, n30509, n30510, n30511,
         n30512, n30513, n30514, n30515, n30516, n30517, n30518, n30519,
         n30520, n30521, n30522, n30523, n30524, n30525, n30526, n30527,
         n30528, n30529, n30530, n30531, n30532, n30533, n30534, n30535,
         n30536, n30537, n30538, n30539, n30540, n30541, n30542, n30543,
         n30544, n30545, n30546, n30547, n30548, n30549, n30550, n30551,
         n30552, n30553, n30554, n30555, n30556, n30557, n30558, n30559,
         n30560, n30561, n30562, n30563, n30564, n30565, n30566, n30567,
         n30568, n30569, n30570, n30571, n30572, n30573, n30574, n30575,
         n30576, n30577, n30578, n30579, n30580, n30581, n30582, n30583,
         n30584, n30585, n30586, n30587, n30588, n30589, n30590, n30591,
         n30592, n30593, n30594, n30595, n30596, n30597, n30598, n30599,
         n30600, n30601, n30602, n30603, n30604, n30605, n30606, n30607,
         n30608, n30609, n30610, n30611, n30612, n30613, n30614, n30615,
         n30616, n30617, n30618, n30619, n30620, n30621, n30622, n30623,
         n30624, n30625, n30626, n30627, n30628, n30629, n30630, n30631,
         n30632, n30633, n30634, n30635, n30636, n30637, n30638, n30639,
         n30640, n30641, n30642, n30643, n30644, n30645, n30646, n30647,
         n30648, n30649, n30650, n30651, n30652, n30653, n30654, n30655,
         n30656, n30657, n30658, n30659, n30660, n30661, n30662, n30663,
         n30664, n30665, n30666, n30667, n30668, n30669, n30670, n30671,
         n30672, n30673, n30674, n30675, n30676, n30677, n30678, n30679,
         n30680, n30681, n30682, n30683, n30684, n30685, n30686, n30687,
         n30688, n30689, n30690, n30691, n30692, n30693, n30694, n30695,
         n30696, n30697, n30698, n30699, n30700, n30701, n30702, n30703,
         n30704, n30705, n30706, n30707, n30708, n30709, n30710, n30711,
         n30712, n30713, n30714, n30715, n30716, n30717, n30718, n30719,
         n30720, n30721, n30722, n30723, n30724, n30725, n30726, n30727,
         n30728, n30729, n30730, n30731, n30732, n30733, n30734, n30735,
         n30736, n30737, n30738, n30739, n30740, n30741, n30742, n30743,
         n30744, n30745, n30746, n30747, n30748, n30749, n30750, n30751,
         n30752, n30753, n30754, n30755, n30756, n30757, n30758, n30759,
         n30760, n30761, n30762, n30763, n30764, n30765, n30766, n30767,
         n30768, n30769, n30770, n30771, n30772, n30773, n30774, n30775,
         n30776, n30777, n30778, n30779, n30780, n30781, n30782, n30783,
         n30784, n30785, n30786, n30787, n30788, n30789, n30790, n30791,
         n30792, n30793, n30794, n30795, n30796, n30797, n30798, n30799,
         n30800, n30801, n30802, n30803, n30804, n30805, n30806, n30807,
         n30808, n30809, n30810, n30811, n30812, n30813, n30814, n30815,
         n30816, n30817, n30818, n30819, n30820, n30821, n30822, n30823,
         n30824, n30825, n30826, n30827, n30828, n30829, n30830, n30831,
         n30832, n30833, n30834, n30835, n30836, n30837, n30838, n30839,
         n30840, n30841, n30842, n30843, n30844, n30845, n30846, n30847,
         n30848, n30849, n30850, n30851, n30852, n30853, n30854, n30855,
         n30856, n30857, n30858, n30859, n30860, n30861, n30862, n30863,
         n30864, n30865, n30866, n30867, n30868, n30869, n30870, n30871,
         n30872, n30873, n30874, n30875, n30876, n30877, n30878, n30879,
         n30880, n30881, n30882, n30883, n30884, n30885, n30886, n30887,
         n30888, n30889, n30890, n30891, n30892, n30893, n30894, n30895,
         n30896, n30897, n30898, n30899, n30900, n30901, n30902, n30903,
         n30904, n30905, n30906, n30907, n30908, n30909, n30910, n30911,
         n30912, n30913, n30914, n30915, n30916, n30917, n30918, n30919,
         n30920, n30921, n30922, n30923, n30924, n30925, n30926, n30927,
         n30928, n30929, n30930, n30931, n30932, n30933, n30934, n30935,
         n30936, n30937, n30938, n30939, n30940, n30941, n30942, n30943,
         n30944, n30945, n30946, n30947, n30948, n30949, n30950, n30951,
         n30952, n30953, n30954, n30955, n30956, n30957, n30958, n30959,
         n30960, n30961, n30962, n30963, n30964, n30965, n30966, n30967,
         n30968, n30969, n30970, n30971, n30972, n30973, n30974, n30975,
         n30976, n30977, n30978, n30979, n30980, n30981, n30982, n30983,
         n30984, n30985, n30986, n30987, n30988, n30989, n30990, n30991,
         n30992, n30993, n30994, n30995, n30996, n30997, n30998, n30999,
         n31000, n31001, n31002, n31003, n31004, n31005, n31006, n31007,
         n31008, n31009, n31010, n31011, n31012, n31013, n31014, n31015,
         n31016, n31017, n31018, n31019, n31020, n31021, n31022, n31023,
         n31024, n31025, n31026, n31027, n31028, n31029, n31030, n31031,
         n31032, n31033, n31034, n31035, n31036, n31037, n31038, n31039,
         n31040, n31041, n31042, n31043, n31044, n31045, n31046, n31047,
         n31048, n31049, n31050, n31051, n31052, n31053, n31054, n31055,
         n31056, n31057, n31058, n31059, n31060, n31061, n31062, n31063,
         n31064, n31065, n31066, n31067, n31068, n31069, n31070, n31071,
         n31072, n31073, n31074, n31075, n31076, n31077, n31078, n31079,
         n31080, n31081, n31082, n31083, n31084, n31085, n31086, n31087,
         n31088, n31089, n31090, n31091, n31092, n31093, n31094, n31095,
         n31096, n31097, n31098, n31099, n31100, n31101, n31102, n31103,
         n31104, n31105, n31106, n31107, n31108, n31109, n31110, n31111,
         n31112, n31113, n31114, n31115, n31116, n31117, n31118, n31119,
         n31120, n31121, n31122, n31123, n31124, n31125, n31126, n31127,
         n31128, n31129, n31130, n31131, n31132, n31133, n31134, n31135,
         n31136, n31137, n31138, n31139, n31140, n31141, n31142, n31143,
         n31144, n31145, n31146, n31147, n31148, n31149, n31150, n31151,
         n31152, n31153, n31154, n31155, n31156, n31157, n31158, n31159,
         n31160, n31161, n31162, n31163, n31164, n31165, n31166, n31167,
         n31168, n31169, n31170, n31171, n31172, n31173, n31174, n31175,
         n31176, n31177, n31178, n31179, n31180, n31181, n31182, n31183,
         n31184, n31185, n31186, n31187, n31188, n31189, n31190, n31191,
         n31192, n31193, n31194, n31195, n31196, n31197, n31198, n31199,
         n31200, n31201, n31202, n31203, n31204, n31205, n31206, n31207,
         n31208, n31209, n31210, n31211, n31212, n31213, n31214, n31215,
         n31216, n31217, n31218, n31219, n31220, n31221, n31222, n31223,
         n31224, n31225, n31226, n31227, n31228, n31229, n31230, n31231,
         n31232, n31233, n31234, n31235, n31236, n31237, n31238, n31239,
         n31240, n31241, n31242, n31243, n31244, n31245, n31246, n31247,
         n31248, n31249, n31250, n31251, n31252, n31253, n31254, n31255,
         n31256, n31257, n31258, n31259, n31260, n31261, n31262, n31263,
         n31264, n31265, n31266, n31267, n31268, n31269, n31270, n31271,
         n31272, n31273, n31274, n31275, n31276, n31277, n31278, n31279,
         n31280, n31281, n31282, n31283, n31284, n31285, n31286, n31287,
         n31288, n31289, n31290, n31291, n31292, n31293, n31294, n31295,
         n31296, n31297, n31298, n31299, n31300, n31301, n31302, n31303,
         n31304, n31305, n31306, n31307, n31308, n31309, n31310, n31311,
         n31312, n31313, n31314, n31315, n31316, n31317, n31318, n31319,
         n31320, n31321, n31322, n31323, n31324, n31325, n31326, n31327,
         n31328, n31329, n31330, n31331, n31332, n31333, n31334, n31335,
         n31336, n31337, n31338, n31339, n31340, n31341, n31342, n31343,
         n31344, n31345, n31346, n31347, n31348, n31349, n31350, n31351,
         n31352, n31353, n31354, n31355, n31356, n31357, n31358, n31359,
         n31360, n31361, n31362, n31363, n31364, n31365, n31366, n31367,
         n31368, n31369, n31370, n31371, n31372, n31373, n31374, n31375,
         n31376, n31377, n31378, n31379, n31380, n31381, n31382, n31383,
         n31384, n31385, n31386, n31387, n31388, n31389, n31390, n31391,
         n31392, n31393, n31394, n31395, n31396, n31397, n31398, n31399,
         n31400, n31401, n31402, n31403, n31404, n31405, n31406, n31407,
         n31408, n31409, n31410, n31411, n31412, n31413, n31414, n31415,
         n31416, n31417, n31418, n31419, n31420, n31421, n31422, n31423,
         n31424, n31425, n31426, n31427, n31428, n31429, n31430, n31431,
         n31432, n31433, n31434, n31435, n31436, n31437, n31438, n31439,
         n31440, n31441, n31442, n31443, n31444, n31445, n31446, n31447,
         n31448, n31449, n31450, n31451, n31452, n31453, n31454, n31455,
         n31456, n31457, n31458, n31459, n31460, n31461, n31462, n31463,
         n31464, n31465, n31466, n31467, n31468, n31469, n31470, n31471,
         n31472, n31473, n31474, n31475, n31476, n31477, n31478, n31479,
         n31480, n31481, n31482, n31483, n31484, n31485, n31486, n31487,
         n31488, n31489, n31490, n31491, n31492, n31493, n31494, n31495,
         n31496, n31497, n31498, n31499, n31500, n31501, n31502, n31503,
         n31504, n31505, n31506, n31507, n31508, n31509, n31510, n31511,
         n31512, n31513, n31514, n31515, n31516, n31517, n31518, n31519,
         n31520, n31521, n31522, n31523, n31524, n31525, n31526, n31527,
         n31528, n31529, n31530, n31531, n31532, n31533, n31534, n31535,
         n31536, n31537, n31538, n31539, n31540, n31541, n31542, n31543,
         n31544, n31545, n31546, n31547, n31548, n31549, n31550, n31551,
         n31552, n31553, n31554, n31555, n31556, n31557, n31558, n31559,
         n31560, n31561, n31562, n31563, n31564, n31565, n31566, n31567,
         n31568, n31569, n31570, n31571, n31572, n31573, n31574, n31575,
         n31576, n31577, n31578, n31579, n31580, n31581, n31582, n31583,
         n31584, n31585, n31586, n31587, n31588, n31589, n31590, n31591,
         n31592, n31593, n31594, n31595, n31596, n31597, n31598, n31599,
         n31600, n31601, n31602, n31603, n31604, n31605, n31606, n31607,
         n31608, n31609, n31610, n31611, n31612, n31613, n31614, n31615,
         n31616, n31617, n31618, n31619, n31620, n31621, n31622, n31623,
         n31624, n31625, n31626, n31627, n31628, n31629, n31630, n31631,
         n31632, n31633, n31634, n31635, n31636, n31637, n31638, n31639,
         n31640, n31641, n31642, n31643, n31644, n31645, n31646, n31647,
         n31648, n31649, n31650, n31651, n31652, n31653, n31654, n31655,
         n31656, n31657, n31658, n31659, n31660, n31661, n31662, n31663,
         n31664, n31665, n31666, n31667, n31668, n31669, n31670, n31671,
         n31672, n31673, n31674, n31675, n31676, n31677, n31678, n31679,
         n31680, n31681, n31682, n31683, n31684, n31685, n31686, n31687,
         n31688, n31689, n31690, n31691, n31692, n31693, n31694, n31695,
         n31696, n31697, n31698, n31699, n31700, n31701, n31702, n31703,
         n31704, n31705, n31706, n31707, n31708, n31709, n31710, n31711,
         n31712, n31713, n31714, n31715, n31716, n31717, n31718, n31719,
         n31720, n31721, n31722, n31723, n31724, n31725, n31726, n31727,
         n31728, n31729, n31730, n31731, n31732, n31733, n31734, n31735,
         n31736, n31737, n31738, n31739, n31740, n31741, n31742, n31743,
         n31744, n31745, n31746, n31747, n31748, n31749, n31750, n31751,
         n31752, n31753, n31754, n31755, n31756, n31757, n31758, n31759,
         n31760, n31761, n31762, n31763, n31764, n31765, n31766, n31767,
         n31768, n31769, n31770, n31771, n31772, n31773, n31774, n31775,
         n31776, n31777, n31778, n31779, n31780, n31781, n31782, n31783,
         n31784, n31785, n31786, n31787, n31788, n31789, n31790, n31791,
         n31792, n31793, n31794, n31795, n31796, n31797, n31798, n31799,
         n31800, n31801, n31802, n31803, n31804, n31805, n31806, n31807,
         n31808, n31809, n31810, n31811, n31812, n31813, n31814, n31815,
         n31816, n31817, n31818, n31819, n31820, n31821, n31822, n31823,
         n31824, n31825, n31826, n31827, n31828, n31829, n31830, n31831,
         n31832, n31833, n31834, n31835, n31836, n31837, n31838, n31839,
         n31840, n31841, n31842, n31843, n31844, n31845, n31846, n31847,
         n31848, n31849, n31850, n31851, n31852, n31853, n31854, n31855,
         n31856, n31857, n31858, n31859, n31860, n31861, n31862, n31863,
         n31864, n31865, n31866, n31867, n31868, n31869, n31870, n31871,
         n31872, n31873, n31874, n31875, n31876, n31877, n31878, n31879,
         n31880, n31881, n31882, n31883, n31884, n31885, n31886, n31887,
         n31888, n31889, n31890, n31891, n31892, n31893, n31894, n31895,
         n31896, n31897, n31898, n31899, n31900, n31901, n31902, n31903,
         n31904, n31905, n31906, n31907, n31908, n31909, n31910, n31911,
         n31912, n31913, n31914, n31915, n31916, n31917, n31918, n31919,
         n31920, n31921, n31922, n31923, n31924, n31925, n31926, n31927,
         n31928, n31929, n31930, n31931, n31932, n31933, n31934, n31935,
         n31936, n31937, n31938, n31939, n31940, n31941, n31942, n31943,
         n31944, n31945, n31946, n31947, n31948, n31949, n31950, n31951,
         n31952, n31953, n31954, n31955, n31956, n31957, n31958, n31959,
         n31960, n31961, n31962, n31963, n31964, n31965, n31966, n31967,
         n31968, n31969, n31970, n31971, n31972, n31973, n31974, n31975,
         n31976, n31977, n31978, n31979, n31980, n31981, n31982, n31983,
         n31984, n31985, n31986, n31987, n31988, n31989, n31990, n31991,
         n31992, n31993, n31994, n31995, n31996, n31997;
  wire   [2:0] c_s;
  wire   [7:0] addr;
  wire   [23:0] act;
  wire   [8:0] cal_cnt;
  wire   [2:0] act_ptr;
  wire   [3:0] set_cnt;
  wire   [1:0] in_cnt;
  wire   [5:0] img_size;
  wire   [3:0] row;
  wire   [3:0] col;
  wire   [3:0] i_row;
  wire   [3:0] i_col;
  wire   [4:0] out_cnt;
  wire   [71:0] template_store;
  wire   [255:0] A67_shift;
  wire   [2047:0] img;
  wire   [7:0] gray_max_out;
  wire   [7:0] gray_avg_out;
  wire   [7:0] gray_weight_out;
  wire   [2:0] act_cnt;
  wire   [3:0] temp_cnt;
  wire   [23:0] rgb_value;
  wire   [7:0] gray_max;
  wire   [7:0] gray_avg;
  wire   [6:0] gray_weight;
  wire   [5:2] img_size_hold;
  wire   [143:0] PE_mul;
  wire   [7:0] m0_DO_reg;
  wire   [7:0] m2_DO_reg;
  wire   [7:0] m1_DO_reg;

  MEM_gray_max m0_U0 ( .A0(addr[0]), .A1(addr[1]), .A2(addr[2]), .A3(addr[3]), 
        .A4(addr[4]), .A5(addr[5]), .A6(addr[6]), .A7(addr[7]), .CK(clk), .CS(
        n11230), .DI0(gray_max[0]), .DI1(gray_max[1]), .DI2(gray_max[2]), 
        .DI3(gray_max[3]), .DI4(gray_max[4]), .DI5(gray_max[5]), .DI6(
        gray_max[6]), .DI7(gray_max[7]), .OE(n11230), .WEB(N25894), .DO0(
        m0_DO_reg[0]), .DO1(m0_DO_reg[1]), .DO2(m0_DO_reg[2]), .DO3(
        m0_DO_reg[3]), .DO4(m0_DO_reg[4]), .DO5(m0_DO_reg[5]), .DO6(
        m0_DO_reg[6]), .DO7(m0_DO_reg[7]) );
  MEM_gray_max m2_U0 ( .A0(addr[0]), .A1(addr[1]), .A2(addr[2]), .A3(addr[3]), 
        .A4(addr[4]), .A5(addr[5]), .A6(addr[6]), .A7(addr[7]), .CK(clk), .CS(
        n11230), .DI0(gray_weight[0]), .DI1(gray_weight[1]), .DI2(
        gray_weight[2]), .DI3(gray_weight[3]), .DI4(gray_weight[4]), .DI5(
        gray_weight[5]), .DI6(gray_weight[6]), .DI7(intadd_8_n1), .OE(n11230), 
        .WEB(N25894), .DO0(m2_DO_reg[0]), .DO1(m2_DO_reg[1]), .DO2(
        m2_DO_reg[2]), .DO3(m2_DO_reg[3]), .DO4(m2_DO_reg[4]), .DO5(
        m2_DO_reg[5]), .DO6(m2_DO_reg[6]), .DO7(m2_DO_reg[7]) );
  MEM_gray_max m1_U0 ( .A0(addr[0]), .A1(addr[1]), .A2(addr[2]), .A3(addr[3]), 
        .A4(addr[4]), .A5(addr[5]), .A6(addr[6]), .A7(addr[7]), .CK(clk), .CS(
        n11230), .DI0(gray_avg[0]), .DI1(gray_avg[1]), .DI2(gray_avg[2]), 
        .DI3(gray_avg[3]), .DI4(gray_avg[4]), .DI5(gray_avg[5]), .DI6(
        gray_avg[6]), .DI7(gray_avg[7]), .OE(n11230), .WEB(N25894), .DO0(
        m1_DO_reg[0]), .DO1(m1_DO_reg[1]), .DO2(m1_DO_reg[2]), .DO3(
        m1_DO_reg[3]), .DO4(m1_DO_reg[4]), .DO5(m1_DO_reg[5]), .DO6(
        m1_DO_reg[6]), .DO7(m1_DO_reg[7]) );
  QDFFRBS in_cnt_reg_0_ ( .D(N25777), .CK(clk), .RB(n13805), .Q(in_cnt[0]) );
  QDFFRBS in_cnt_reg_1_ ( .D(N25778), .CK(clk), .RB(n13805), .Q(in_cnt[1]) );
  QDFFRBS img_size_reg_5_ ( .D(n13639), .CK(clk), .RB(n13805), .Q(img_size[5])
         );
  QDFFRBS c_s_reg_2_ ( .D(n30029), .CK(clk), .RB(n13805), .Q(c_s[2]) );
  QDFFRBS c_s_reg_1_ ( .D(n30027), .CK(clk), .RB(n13805), .Q(c_s[1]) );
  QDFFRBS out_cnt_reg_2_ ( .D(n13680), .CK(clk), .RB(n13805), .Q(out_cnt[2])
         );
  QDFFRBS out_cnt_reg_3_ ( .D(n13679), .CK(clk), .RB(n13805), .Q(out_cnt[3])
         );
  QDFFRBS addr_reg_7_ ( .D(n13633), .CK(clk), .RB(n13805), .Q(addr[7]) );
  QDFFRBS addr_reg_0_ ( .D(n13632), .CK(clk), .RB(n13805), .Q(addr[0]) );
  QDFFRBS addr_reg_1_ ( .D(n13631), .CK(clk), .RB(n13805), .Q(addr[1]) );
  QDFFRBS addr_reg_2_ ( .D(n13630), .CK(clk), .RB(n13805), .Q(addr[2]) );
  QDFFRBS addr_reg_4_ ( .D(n13628), .CK(clk), .RB(n13805), .Q(addr[4]) );
  QDFFRBS addr_reg_5_ ( .D(n13627), .CK(clk), .RB(n13805), .Q(addr[5]) );
  QDFFRBS cal_cnt_reg_1_ ( .D(n13654), .CK(clk), .RB(n13805), .Q(cal_cnt[1])
         );
  QDFFRBS cal_cnt_reg_0_ ( .D(n13653), .CK(clk), .RB(n13805), .Q(cal_cnt[0])
         );
  QDFFRBS cal_cnt_reg_2_ ( .D(n13652), .CK(clk), .RB(n13805), .Q(cal_cnt[2])
         );
  QDFFRBS cal_cnt_reg_3_ ( .D(n13651), .CK(clk), .RB(n13805), .Q(cal_cnt[3])
         );
  QDFFRBS cal_cnt_reg_4_ ( .D(n13650), .CK(clk), .RB(n13805), .Q(cal_cnt[4])
         );
  QDFFRBS cal_cnt_reg_5_ ( .D(n13649), .CK(clk), .RB(n13805), .Q(cal_cnt[5])
         );
  QDFFRBS cal_cnt_reg_6_ ( .D(n13648), .CK(clk), .RB(n13805), .Q(cal_cnt[6])
         );
  QDFFRBS cal_cnt_reg_7_ ( .D(n13647), .CK(clk), .RB(n13805), .Q(cal_cnt[7])
         );
  QDFFRBS cal_cnt_reg_8_ ( .D(n13646), .CK(clk), .RB(n13805), .Q(cal_cnt[8])
         );
  QDFFRBS set_cnt_reg_0_ ( .D(n13940), .CK(clk), .RB(n13805), .Q(set_cnt[0])
         );
  QDFFRBS set_cnt_reg_1_ ( .D(n13636), .CK(clk), .RB(n13805), .Q(set_cnt[1])
         );
  QDFFRBS set_cnt_reg_2_ ( .D(n13635), .CK(clk), .RB(n13805), .Q(set_cnt[2])
         );
  QDFFRBS set_cnt_reg_3_ ( .D(n13634), .CK(clk), .RB(n13805), .Q(set_cnt[3])
         );
  QDFFRBS temp_cnt_reg_0_ ( .D(n13625), .CK(clk), .RB(n13805), .Q(temp_cnt[0])
         );
  QDFFRBS temp_cnt_reg_2_ ( .D(n13623), .CK(clk), .RB(n13805), .Q(temp_cnt[2])
         );
  QDFFRBS temp_cnt_reg_3_ ( .D(n13622), .CK(clk), .RB(n13805), .Q(temp_cnt[3])
         );
  QDFFRBS act_cnt_reg_0_ ( .D(n13688), .CK(clk), .RB(n13805), .Q(act_cnt[0])
         );
  QDFFRBS act_cnt_reg_1_ ( .D(n13687), .CK(clk), .RB(n13805), .Q(act_cnt[1])
         );
  QDFFRBS act_cnt_reg_2_ ( .D(n13686), .CK(clk), .RB(n13805), .Q(act_cnt[2])
         );
  QDFFRBS act_reg_7__0_ ( .D(n13678), .CK(clk), .RB(n13805), .Q(act[0]) );
  QDFFRBS act_reg_7__2_ ( .D(n13677), .CK(clk), .RB(n13805), .Q(act[2]) );
  QDFFRBS act_reg_7__1_ ( .D(n13676), .CK(clk), .RB(n30035), .Q(act[1]) );
  QDFFRBS act_reg_6__0_ ( .D(n13675), .CK(clk), .RB(n13805), .Q(act[3]) );
  QDFFRBS act_reg_6__2_ ( .D(n13674), .CK(clk), .RB(n13805), .Q(act[5]) );
  QDFFRBS act_reg_6__1_ ( .D(n13673), .CK(clk), .RB(n13805), .Q(act[4]) );
  QDFFRBS act_reg_5__0_ ( .D(n13672), .CK(clk), .RB(n13805), .Q(act[6]) );
  QDFFRBS act_reg_5__2_ ( .D(n13671), .CK(clk), .RB(n13805), .Q(act[8]) );
  QDFFRBS act_reg_5__1_ ( .D(n13670), .CK(clk), .RB(n13805), .Q(act[7]) );
  QDFFRBS act_reg_4__0_ ( .D(n13669), .CK(clk), .RB(n13805), .Q(act[9]) );
  QDFFRBS act_reg_4__2_ ( .D(n13668), .CK(clk), .RB(n13805), .Q(act[11]) );
  QDFFRBS act_reg_4__1_ ( .D(n13667), .CK(clk), .RB(n13805), .Q(act[10]) );
  QDFFRBS act_reg_3__0_ ( .D(n13666), .CK(clk), .RB(n13805), .Q(act[12]) );
  QDFFRBS act_reg_3__2_ ( .D(n13665), .CK(clk), .RB(n13805), .Q(act[14]) );
  QDFFRBS act_reg_3__1_ ( .D(n13664), .CK(clk), .RB(n13805), .Q(act[13]) );
  QDFFRBS act_reg_2__0_ ( .D(n13663), .CK(clk), .RB(n13805), .Q(act[15]) );
  QDFFRBS act_reg_2__2_ ( .D(n13662), .CK(clk), .RB(n13805), .Q(act[17]) );
  QDFFRBS act_reg_2__1_ ( .D(n13661), .CK(clk), .RB(n13805), .Q(act[16]) );
  QDFFRBS act_reg_1__0_ ( .D(n13660), .CK(clk), .RB(n13805), .Q(act[18]) );
  QDFFRBS act_reg_1__2_ ( .D(n13659), .CK(clk), .RB(n13805), .Q(act[20]) );
  QDFFRBS act_reg_1__1_ ( .D(n13658), .CK(clk), .RB(n13805), .Q(act[19]) );
  QDFFRBS act_reg_0__0_ ( .D(n13657), .CK(clk), .RB(n13805), .Q(act[21]) );
  QDFFRBS act_reg_0__2_ ( .D(n13656), .CK(clk), .RB(n13805), .Q(act[23]) );
  QDFFRBS act_reg_0__1_ ( .D(n13655), .CK(clk), .RB(n13805), .Q(act[22]) );
  QDFFRBS act_ptr_reg_1_ ( .D(n13645), .CK(clk), .RB(n13805), .Q(act_ptr[1])
         );
  QDFFRBS act_ptr_reg_2_ ( .D(n13684), .CK(clk), .RB(n13805), .Q(act_ptr[2])
         );
  QDFFRBS row_reg_0_ ( .D(n13619), .CK(clk), .RB(n13805), .Q(row[0]) );
  QDFFRBS row_reg_1_ ( .D(n13616), .CK(clk), .RB(n13805), .Q(row[1]) );
  QDFFRBS row_reg_2_ ( .D(n13617), .CK(clk), .RB(n13805), .Q(row[2]) );
  QDFFRBS row_reg_3_ ( .D(n13618), .CK(clk), .RB(n13805), .Q(row[3]) );
  QDFFRBS col_reg_0_ ( .D(n13615), .CK(clk), .RB(n13805), .Q(col[0]) );
  QDFFRBS col_reg_2_ ( .D(n13614), .CK(clk), .RB(n13805), .Q(col[2]) );
  QDFFRBS col_reg_3_ ( .D(n13620), .CK(clk), .RB(n13805), .Q(col[3]) );
  QDFFRBS template_store_reg_0__7_ ( .D(n13605), .CK(clk), .RB(n13805), .Q(
        template_store[71]) );
  QDFFRBS template_store_reg_0__6_ ( .D(n13604), .CK(clk), .RB(n13805), .Q(
        template_store[70]) );
  QDFFRBS template_store_reg_0__5_ ( .D(n13603), .CK(clk), .RB(n13805), .Q(
        template_store[69]) );
  QDFFRBS template_store_reg_0__4_ ( .D(n13602), .CK(clk), .RB(n13805), .Q(
        template_store[68]) );
  QDFFRBS template_store_reg_0__3_ ( .D(n13601), .CK(clk), .RB(n13805), .Q(
        template_store[67]) );
  QDFFRBS template_store_reg_0__2_ ( .D(n13600), .CK(clk), .RB(rst_n), .Q(
        template_store[66]) );
  QDFFRBS template_store_reg_0__1_ ( .D(n13599), .CK(clk), .RB(rst_n), .Q(
        template_store[65]) );
  QDFFRBS template_store_reg_0__0_ ( .D(n13598), .CK(clk), .RB(rst_n), .Q(
        template_store[64]) );
  QDFFRBS template_store_reg_1__7_ ( .D(n13597), .CK(clk), .RB(rst_n), .Q(
        template_store[63]) );
  QDFFRBS template_store_reg_1__6_ ( .D(n13596), .CK(clk), .RB(rst_n), .Q(
        template_store[62]) );
  QDFFRBS template_store_reg_1__5_ ( .D(n13595), .CK(clk), .RB(n13805), .Q(
        template_store[61]) );
  QDFFRBS template_store_reg_1__4_ ( .D(n13594), .CK(clk), .RB(n13805), .Q(
        template_store[60]) );
  QDFFRBS template_store_reg_1__3_ ( .D(n13593), .CK(clk), .RB(n13805), .Q(
        template_store[59]) );
  QDFFRBS template_store_reg_1__2_ ( .D(n13592), .CK(clk), .RB(n30035), .Q(
        template_store[58]) );
  QDFFRBS template_store_reg_1__1_ ( .D(n13591), .CK(clk), .RB(n13805), .Q(
        template_store[57]) );
  QDFFRBS template_store_reg_1__0_ ( .D(n13590), .CK(clk), .RB(n30034), .Q(
        template_store[56]) );
  QDFFRBS template_store_reg_2__7_ ( .D(n13589), .CK(clk), .RB(n30034), .Q(
        template_store[55]) );
  QDFFRBS template_store_reg_2__6_ ( .D(n13588), .CK(clk), .RB(n30034), .Q(
        template_store[54]) );
  QDFFRBS template_store_reg_2__5_ ( .D(n13587), .CK(clk), .RB(n30034), .Q(
        template_store[53]) );
  QDFFRBS template_store_reg_2__4_ ( .D(n13586), .CK(clk), .RB(n30034), .Q(
        template_store[52]) );
  QDFFRBS template_store_reg_2__3_ ( .D(n13585), .CK(clk), .RB(n30034), .Q(
        template_store[51]) );
  QDFFRBS template_store_reg_2__2_ ( .D(n13584), .CK(clk), .RB(n30034), .Q(
        template_store[50]) );
  QDFFRBS template_store_reg_2__1_ ( .D(n13583), .CK(clk), .RB(n30034), .Q(
        template_store[49]) );
  QDFFRBS template_store_reg_2__0_ ( .D(n13582), .CK(clk), .RB(n30034), .Q(
        template_store[48]) );
  QDFFRBS template_store_reg_3__7_ ( .D(n13581), .CK(clk), .RB(n30034), .Q(
        template_store[47]) );
  QDFFRBS template_store_reg_3__6_ ( .D(n13580), .CK(clk), .RB(n13805), .Q(
        template_store[46]) );
  QDFFRBS template_store_reg_3__5_ ( .D(n13579), .CK(clk), .RB(n13805), .Q(
        template_store[45]) );
  QDFFRBS template_store_reg_3__4_ ( .D(n13578), .CK(clk), .RB(n13805), .Q(
        template_store[44]) );
  QDFFRBS template_store_reg_3__3_ ( .D(n13577), .CK(clk), .RB(n13805), .Q(
        template_store[43]) );
  QDFFRBS template_store_reg_3__2_ ( .D(n13576), .CK(clk), .RB(n13805), .Q(
        template_store[42]) );
  QDFFRBS template_store_reg_3__1_ ( .D(n13575), .CK(clk), .RB(n13805), .Q(
        template_store[41]) );
  QDFFRBS template_store_reg_3__0_ ( .D(n13574), .CK(clk), .RB(n13805), .Q(
        template_store[40]) );
  QDFFRBS template_store_reg_4__7_ ( .D(n13573), .CK(clk), .RB(n13805), .Q(
        template_store[39]) );
  QDFFRBS template_store_reg_4__6_ ( .D(n13572), .CK(clk), .RB(n13805), .Q(
        template_store[38]) );
  QDFFRBS template_store_reg_4__5_ ( .D(n13571), .CK(clk), .RB(n13805), .Q(
        template_store[37]) );
  QDFFRBS template_store_reg_4__4_ ( .D(n13570), .CK(clk), .RB(n13805), .Q(
        template_store[36]) );
  QDFFRBS template_store_reg_4__3_ ( .D(n13569), .CK(clk), .RB(n13805), .Q(
        template_store[35]) );
  QDFFRBS template_store_reg_4__2_ ( .D(n13568), .CK(clk), .RB(n13805), .Q(
        template_store[34]) );
  QDFFRBS template_store_reg_4__1_ ( .D(n13567), .CK(clk), .RB(n13805), .Q(
        template_store[33]) );
  QDFFRBS template_store_reg_4__0_ ( .D(n13566), .CK(clk), .RB(n13805), .Q(
        template_store[32]) );
  QDFFRBS template_store_reg_5__7_ ( .D(n13565), .CK(clk), .RB(n13805), .Q(
        template_store[31]) );
  QDFFRBS template_store_reg_5__6_ ( .D(n13564), .CK(clk), .RB(n13805), .Q(
        template_store[30]) );
  QDFFRBS template_store_reg_5__5_ ( .D(n13563), .CK(clk), .RB(n13805), .Q(
        template_store[29]) );
  QDFFRBS template_store_reg_5__4_ ( .D(n13562), .CK(clk), .RB(n13805), .Q(
        template_store[28]) );
  QDFFRBS template_store_reg_5__3_ ( .D(n13561), .CK(clk), .RB(n13805), .Q(
        template_store[27]) );
  QDFFRBS template_store_reg_5__2_ ( .D(n13560), .CK(clk), .RB(n13805), .Q(
        template_store[26]) );
  QDFFRBS template_store_reg_5__1_ ( .D(n13559), .CK(clk), .RB(n13805), .Q(
        template_store[25]) );
  QDFFRBS template_store_reg_5__0_ ( .D(n13558), .CK(clk), .RB(n13805), .Q(
        template_store[24]) );
  QDFFRBS template_store_reg_6__7_ ( .D(n13557), .CK(clk), .RB(n13805), .Q(
        template_store[23]) );
  QDFFRBS template_store_reg_6__6_ ( .D(n13556), .CK(clk), .RB(n13805), .Q(
        template_store[22]) );
  QDFFRBS template_store_reg_6__5_ ( .D(n13555), .CK(clk), .RB(n13805), .Q(
        template_store[21]) );
  QDFFRBS template_store_reg_6__4_ ( .D(n13554), .CK(clk), .RB(n13805), .Q(
        template_store[20]) );
  QDFFRBS template_store_reg_6__3_ ( .D(n13553), .CK(clk), .RB(n13805), .Q(
        template_store[19]) );
  QDFFRBS template_store_reg_6__2_ ( .D(n13552), .CK(clk), .RB(n30034), .Q(
        template_store[18]) );
  QDFFRBS template_store_reg_6__1_ ( .D(n13551), .CK(clk), .RB(n30034), .Q(
        template_store[17]) );
  QDFFRBS template_store_reg_6__0_ ( .D(n13550), .CK(clk), .RB(n30034), .Q(
        template_store[16]) );
  QDFFRBS template_store_reg_7__7_ ( .D(n13549), .CK(clk), .RB(n30034), .Q(
        template_store[15]) );
  QDFFRBS template_store_reg_7__6_ ( .D(n13548), .CK(clk), .RB(n30034), .Q(
        template_store[14]) );
  QDFFRBS template_store_reg_7__5_ ( .D(n13547), .CK(clk), .RB(n30034), .Q(
        template_store[13]) );
  QDFFRBS template_store_reg_7__4_ ( .D(n13546), .CK(clk), .RB(n30034), .Q(
        template_store[12]) );
  QDFFRBS template_store_reg_7__3_ ( .D(n13545), .CK(clk), .RB(n30034), .Q(
        template_store[11]) );
  QDFFRBS template_store_reg_7__2_ ( .D(n13544), .CK(clk), .RB(n30034), .Q(
        template_store[10]) );
  QDFFRBS template_store_reg_7__1_ ( .D(n13543), .CK(clk), .RB(n30034), .Q(
        template_store[9]) );
  QDFFRBS template_store_reg_7__0_ ( .D(n13542), .CK(clk), .RB(n30034), .Q(
        template_store[8]) );
  QDFFRBS template_store_reg_8__7_ ( .D(n13541), .CK(clk), .RB(n30034), .Q(
        template_store[7]) );
  QDFFRBS template_store_reg_8__6_ ( .D(n13540), .CK(clk), .RB(n30034), .Q(
        template_store[6]) );
  QDFFRBS template_store_reg_8__5_ ( .D(n13539), .CK(clk), .RB(n30035), .Q(
        template_store[5]) );
  QDFFRBS template_store_reg_8__4_ ( .D(n13538), .CK(clk), .RB(n30035), .Q(
        template_store[4]) );
  QDFFRBS template_store_reg_8__3_ ( .D(n13537), .CK(clk), .RB(n30035), .Q(
        template_store[3]) );
  QDFFRBS template_store_reg_8__2_ ( .D(n13536), .CK(clk), .RB(n30035), .Q(
        template_store[2]) );
  QDFFRBS template_store_reg_8__1_ ( .D(n13535), .CK(clk), .RB(n30035), .Q(
        template_store[1]) );
  QDFFRBS template_store_reg_8__0_ ( .D(n13534), .CK(clk), .RB(n30035), .Q(
        template_store[0]) );
  QDFFRBS rgb_value_reg_23_ ( .D(n11228), .CK(clk), .RB(n30035), .Q(
        rgb_value[23]) );
  QDFFRBS rgb_value_reg_22_ ( .D(n11227), .CK(clk), .RB(n30035), .Q(
        rgb_value[22]) );
  QDFFRBS rgb_value_reg_21_ ( .D(n11226), .CK(clk), .RB(n30035), .Q(
        rgb_value[21]) );
  QDFFRBS rgb_value_reg_20_ ( .D(n11225), .CK(clk), .RB(n30035), .Q(
        rgb_value[20]) );
  QDFFRBS rgb_value_reg_19_ ( .D(n11224), .CK(clk), .RB(n30035), .Q(
        rgb_value[19]) );
  QDFFRBS rgb_value_reg_18_ ( .D(n11223), .CK(clk), .RB(n30035), .Q(
        rgb_value[18]) );
  QDFFRBS rgb_value_reg_17_ ( .D(n11222), .CK(clk), .RB(n30035), .Q(
        rgb_value[17]) );
  QDFFRBS rgb_value_reg_16_ ( .D(n11221), .CK(clk), .RB(n30035), .Q(
        rgb_value[16]) );
  QDFFRBS rgb_value_reg_13_ ( .D(n11218), .CK(clk), .RB(n30035), .Q(
        rgb_value[13]) );
  QDFFRBS rgb_value_reg_12_ ( .D(n11217), .CK(clk), .RB(n30035), .Q(
        rgb_value[12]) );
  QDFFRBS rgb_value_reg_11_ ( .D(n11216), .CK(clk), .RB(n30035), .Q(
        rgb_value[11]) );
  QDFFRBS rgb_value_reg_10_ ( .D(n11215), .CK(clk), .RB(n30035), .Q(
        rgb_value[10]) );
  QDFFRBS rgb_value_reg_9_ ( .D(n11214), .CK(clk), .RB(n30035), .Q(
        rgb_value[9]) );
  QDFFRBS rgb_value_reg_8_ ( .D(n11213), .CK(clk), .RB(n30035), .Q(
        rgb_value[8]) );
  QDFFRBS rgb_value_reg_5_ ( .D(n11210), .CK(clk), .RB(n30035), .Q(
        rgb_value[5]) );
  QDFFRBS rgb_value_reg_3_ ( .D(n11208), .CK(clk), .RB(rst_n), .Q(rgb_value[3]) );
  QDFFRBS rgb_value_reg_2_ ( .D(n11207), .CK(clk), .RB(n30035), .Q(
        rgb_value[2]) );
  QDFFRBS rgb_value_reg_1_ ( .D(n11206), .CK(clk), .RB(n30035), .Q(
        rgb_value[1]) );
  QDFFRBS rgb_value_reg_0_ ( .D(n11205), .CK(clk), .RB(n30035), .Q(
        rgb_value[0]) );
  QDFFRBS img_size_hold_reg_5_ ( .D(n11204), .CK(clk), .RB(n30035), .Q(
        img_size_hold[5]) );
  QDFFRBS img_size_hold_reg_4_ ( .D(n11203), .CK(clk), .RB(n30035), .Q(
        img_size_hold[4]) );
  QDFFRBS img_size_hold_reg_3_ ( .D(n11202), .CK(clk), .RB(n30035), .Q(
        img_size_hold[3]) );
  QDFFRBS img_size_hold_reg_2_ ( .D(n11201), .CK(clk), .RB(n30035), .Q(
        img_size_hold[2]) );
  QDFFS act_delay1_reg ( .D(n30026), .CK(clk), .Q(act_delay1) );
  QDFFS act_delay2_reg ( .D(act_delay1), .CK(clk), .Q(act_delay2) );
  QDFFS PE_mul_reg_8__0_ ( .D(PE_N128), .CK(clk), .Q(PE_mul[0]) );
  QDFFS PE_mul_reg_8__1_ ( .D(PE_N129), .CK(clk), .Q(PE_mul[1]) );
  QDFFS PE_mul_reg_8__2_ ( .D(PE_N130), .CK(clk), .Q(PE_mul[2]) );
  QDFFS PE_mul_reg_8__3_ ( .D(PE_N131), .CK(clk), .Q(PE_mul[3]) );
  QDFFS PE_mul_reg_8__4_ ( .D(PE_N132), .CK(clk), .Q(PE_mul[4]) );
  QDFFS PE_mul_reg_8__5_ ( .D(PE_N133), .CK(clk), .Q(PE_mul[5]) );
  QDFFS PE_mul_reg_8__6_ ( .D(PE_N134), .CK(clk), .Q(PE_mul[6]) );
  QDFFS PE_mul_reg_8__7_ ( .D(PE_N135), .CK(clk), .Q(PE_mul[7]) );
  QDFFS PE_mul_reg_8__8_ ( .D(PE_N136), .CK(clk), .Q(PE_mul[8]) );
  QDFFS PE_mul_reg_8__9_ ( .D(PE_N137), .CK(clk), .Q(PE_mul[9]) );
  QDFFS PE_mul_reg_8__10_ ( .D(PE_N138), .CK(clk), .Q(PE_mul[10]) );
  QDFFS PE_mul_reg_8__11_ ( .D(PE_N139), .CK(clk), .Q(PE_mul[11]) );
  QDFFS PE_mul_reg_8__12_ ( .D(PE_N140), .CK(clk), .Q(PE_mul[12]) );
  QDFFS PE_mul_reg_8__13_ ( .D(PE_N141), .CK(clk), .Q(PE_mul[13]) );
  QDFFS PE_mul_reg_8__14_ ( .D(PE_N142), .CK(clk), .Q(PE_mul[14]) );
  QDFFS PE_mul_reg_8__15_ ( .D(PE_N143), .CK(clk), .Q(PE_mul[15]) );
  QDFFS PE_mul_reg_7__0_ ( .D(PE_N112), .CK(clk), .Q(PE_mul[16]) );
  QDFFS PE_mul_reg_7__1_ ( .D(PE_N113), .CK(clk), .Q(PE_mul[17]) );
  QDFFS PE_mul_reg_7__2_ ( .D(PE_N114), .CK(clk), .Q(PE_mul[18]) );
  QDFFS PE_mul_reg_7__3_ ( .D(PE_N115), .CK(clk), .Q(PE_mul[19]) );
  QDFFS PE_mul_reg_7__4_ ( .D(PE_N116), .CK(clk), .Q(PE_mul[20]) );
  QDFFS PE_mul_reg_7__5_ ( .D(PE_N117), .CK(clk), .Q(PE_mul[21]) );
  QDFFS PE_mul_reg_7__6_ ( .D(PE_N118), .CK(clk), .Q(PE_mul[22]) );
  QDFFS PE_mul_reg_7__7_ ( .D(PE_N119), .CK(clk), .Q(PE_mul[23]) );
  QDFFS PE_mul_reg_7__8_ ( .D(PE_N120), .CK(clk), .Q(PE_mul[24]) );
  QDFFS PE_mul_reg_7__9_ ( .D(PE_N121), .CK(clk), .Q(PE_mul[25]) );
  QDFFS PE_mul_reg_7__10_ ( .D(PE_N122), .CK(clk), .Q(PE_mul[26]) );
  QDFFS PE_mul_reg_7__11_ ( .D(PE_N123), .CK(clk), .Q(PE_mul[27]) );
  QDFFS PE_mul_reg_7__12_ ( .D(PE_N124), .CK(clk), .Q(PE_mul[28]) );
  QDFFS PE_mul_reg_7__13_ ( .D(PE_N125), .CK(clk), .Q(PE_mul[29]) );
  QDFFS PE_mul_reg_7__14_ ( .D(PE_N126), .CK(clk), .Q(PE_mul[30]) );
  QDFFS PE_mul_reg_7__15_ ( .D(PE_N127), .CK(clk), .Q(PE_mul[31]) );
  QDFFS PE_mul_reg_6__0_ ( .D(PE_N96), .CK(clk), .Q(PE_mul[32]) );
  QDFFS PE_mul_reg_6__1_ ( .D(PE_N97), .CK(clk), .Q(PE_mul[33]) );
  QDFFS PE_mul_reg_6__2_ ( .D(PE_N98), .CK(clk), .Q(PE_mul[34]) );
  QDFFS PE_mul_reg_6__3_ ( .D(PE_N99), .CK(clk), .Q(PE_mul[35]) );
  QDFFS PE_mul_reg_6__4_ ( .D(PE_N100), .CK(clk), .Q(PE_mul[36]) );
  QDFFS PE_mul_reg_6__5_ ( .D(PE_N101), .CK(clk), .Q(PE_mul[37]) );
  QDFFS PE_mul_reg_6__6_ ( .D(PE_N102), .CK(clk), .Q(PE_mul[38]) );
  QDFFS PE_mul_reg_6__7_ ( .D(PE_N103), .CK(clk), .Q(PE_mul[39]) );
  QDFFS PE_mul_reg_6__8_ ( .D(PE_N104), .CK(clk), .Q(PE_mul[40]) );
  QDFFS PE_mul_reg_6__9_ ( .D(PE_N105), .CK(clk), .Q(PE_mul[41]) );
  QDFFS PE_mul_reg_6__10_ ( .D(PE_N106), .CK(clk), .Q(PE_mul[42]) );
  QDFFS PE_mul_reg_6__11_ ( .D(PE_N107), .CK(clk), .Q(PE_mul[43]) );
  QDFFS PE_mul_reg_6__12_ ( .D(PE_N108), .CK(clk), .Q(PE_mul[44]) );
  QDFFS PE_mul_reg_6__13_ ( .D(PE_N109), .CK(clk), .Q(PE_mul[45]) );
  QDFFS PE_mul_reg_6__14_ ( .D(PE_N110), .CK(clk), .Q(PE_mul[46]) );
  QDFFS PE_mul_reg_6__15_ ( .D(PE_N111), .CK(clk), .Q(PE_mul[47]) );
  QDFFS PE_mul_reg_5__0_ ( .D(PE_N80), .CK(clk), .Q(PE_mul[48]) );
  QDFFS PE_mul_reg_5__1_ ( .D(PE_N81), .CK(clk), .Q(PE_mul[49]) );
  QDFFS PE_mul_reg_5__2_ ( .D(PE_N82), .CK(clk), .Q(PE_mul[50]) );
  QDFFS PE_mul_reg_5__3_ ( .D(PE_N83), .CK(clk), .Q(PE_mul[51]) );
  QDFFS PE_mul_reg_5__4_ ( .D(PE_N84), .CK(clk), .Q(PE_mul[52]) );
  QDFFS PE_mul_reg_5__5_ ( .D(PE_N85), .CK(clk), .Q(PE_mul[53]) );
  QDFFS PE_mul_reg_5__6_ ( .D(PE_N86), .CK(clk), .Q(PE_mul[54]) );
  QDFFS PE_mul_reg_5__7_ ( .D(PE_N87), .CK(clk), .Q(PE_mul[55]) );
  QDFFS PE_mul_reg_5__8_ ( .D(PE_N88), .CK(clk), .Q(PE_mul[56]) );
  QDFFS PE_mul_reg_5__9_ ( .D(PE_N89), .CK(clk), .Q(PE_mul[57]) );
  QDFFS PE_mul_reg_5__10_ ( .D(PE_N90), .CK(clk), .Q(PE_mul[58]) );
  QDFFS PE_mul_reg_5__11_ ( .D(PE_N91), .CK(clk), .Q(PE_mul[59]) );
  QDFFS PE_mul_reg_5__12_ ( .D(PE_N92), .CK(clk), .Q(PE_mul[60]) );
  QDFFS PE_mul_reg_5__13_ ( .D(PE_N93), .CK(clk), .Q(PE_mul[61]) );
  QDFFS PE_mul_reg_5__14_ ( .D(PE_N94), .CK(clk), .Q(PE_mul[62]) );
  QDFFS PE_mul_reg_4__0_ ( .D(PE_N64), .CK(clk), .Q(PE_mul[64]) );
  QDFFS PE_mul_reg_4__1_ ( .D(PE_N65), .CK(clk), .Q(PE_mul[65]) );
  QDFFS PE_mul_reg_4__2_ ( .D(PE_N66), .CK(clk), .Q(PE_mul[66]) );
  QDFFS PE_mul_reg_4__3_ ( .D(PE_N67), .CK(clk), .Q(PE_mul[67]) );
  QDFFS PE_mul_reg_4__4_ ( .D(PE_N68), .CK(clk), .Q(PE_mul[68]) );
  QDFFS PE_mul_reg_4__5_ ( .D(PE_N69), .CK(clk), .Q(PE_mul[69]) );
  QDFFS PE_mul_reg_4__6_ ( .D(PE_N70), .CK(clk), .Q(PE_mul[70]) );
  QDFFS PE_mul_reg_4__7_ ( .D(PE_N71), .CK(clk), .Q(PE_mul[71]) );
  QDFFS PE_mul_reg_4__8_ ( .D(PE_N72), .CK(clk), .Q(PE_mul[72]) );
  QDFFS PE_mul_reg_4__9_ ( .D(PE_N73), .CK(clk), .Q(PE_mul[73]) );
  QDFFS PE_mul_reg_4__10_ ( .D(PE_N74), .CK(clk), .Q(PE_mul[74]) );
  QDFFS PE_mul_reg_4__11_ ( .D(PE_N75), .CK(clk), .Q(PE_mul[75]) );
  QDFFS PE_mul_reg_4__12_ ( .D(PE_N76), .CK(clk), .Q(PE_mul[76]) );
  QDFFS PE_mul_reg_4__13_ ( .D(PE_N77), .CK(clk), .Q(PE_mul[77]) );
  QDFFS PE_mul_reg_4__14_ ( .D(PE_N78), .CK(clk), .Q(PE_mul[78]) );
  QDFFS PE_mul_reg_3__0_ ( .D(PE_N48), .CK(clk), .Q(PE_mul[80]) );
  QDFFS PE_mul_reg_3__1_ ( .D(PE_N49), .CK(clk), .Q(PE_mul[81]) );
  QDFFS PE_mul_reg_3__2_ ( .D(PE_N50), .CK(clk), .Q(PE_mul[82]) );
  QDFFS PE_mul_reg_3__3_ ( .D(PE_N51), .CK(clk), .Q(PE_mul[83]) );
  QDFFS PE_mul_reg_3__4_ ( .D(PE_N52), .CK(clk), .Q(PE_mul[84]) );
  QDFFS PE_mul_reg_3__5_ ( .D(PE_N53), .CK(clk), .Q(PE_mul[85]) );
  QDFFS PE_mul_reg_3__6_ ( .D(PE_N54), .CK(clk), .Q(PE_mul[86]) );
  QDFFS PE_mul_reg_3__7_ ( .D(PE_N55), .CK(clk), .Q(PE_mul[87]) );
  QDFFS PE_mul_reg_3__8_ ( .D(PE_N56), .CK(clk), .Q(PE_mul[88]) );
  QDFFS PE_mul_reg_3__9_ ( .D(PE_N57), .CK(clk), .Q(PE_mul[89]) );
  QDFFS PE_mul_reg_3__10_ ( .D(PE_N58), .CK(clk), .Q(PE_mul[90]) );
  QDFFS PE_mul_reg_3__11_ ( .D(PE_N59), .CK(clk), .Q(PE_mul[91]) );
  QDFFS PE_mul_reg_3__12_ ( .D(PE_N60), .CK(clk), .Q(PE_mul[92]) );
  QDFFS PE_mul_reg_3__13_ ( .D(PE_N61), .CK(clk), .Q(PE_mul[93]) );
  QDFFS PE_mul_reg_3__14_ ( .D(PE_N62), .CK(clk), .Q(PE_mul[94]) );
  QDFFS PE_mul_reg_2__0_ ( .D(PE_N32), .CK(clk), .Q(PE_mul[96]) );
  QDFFS PE_mul_reg_2__1_ ( .D(PE_N33), .CK(clk), .Q(PE_mul[97]) );
  QDFFS PE_mul_reg_2__2_ ( .D(PE_N34), .CK(clk), .Q(PE_mul[98]) );
  QDFFS PE_mul_reg_2__3_ ( .D(PE_N35), .CK(clk), .Q(PE_mul[99]) );
  QDFFS PE_mul_reg_2__4_ ( .D(PE_N36), .CK(clk), .Q(PE_mul[100]) );
  QDFFS PE_mul_reg_2__5_ ( .D(PE_N37), .CK(clk), .Q(PE_mul[101]) );
  QDFFS PE_mul_reg_2__6_ ( .D(PE_N38), .CK(clk), .Q(PE_mul[102]) );
  QDFFS PE_mul_reg_2__7_ ( .D(PE_N39), .CK(clk), .Q(PE_mul[103]) );
  QDFFS PE_mul_reg_2__8_ ( .D(PE_N40), .CK(clk), .Q(PE_mul[104]) );
  QDFFS PE_mul_reg_2__9_ ( .D(PE_N41), .CK(clk), .Q(PE_mul[105]) );
  QDFFS PE_mul_reg_2__10_ ( .D(PE_N42), .CK(clk), .Q(PE_mul[106]) );
  QDFFS PE_mul_reg_2__11_ ( .D(PE_N43), .CK(clk), .Q(PE_mul[107]) );
  QDFFS PE_mul_reg_2__12_ ( .D(PE_N44), .CK(clk), .Q(PE_mul[108]) );
  QDFFS PE_mul_reg_2__13_ ( .D(PE_N45), .CK(clk), .Q(PE_mul[109]) );
  QDFFS PE_mul_reg_2__14_ ( .D(PE_N46), .CK(clk), .Q(PE_mul[110]) );
  QDFFS PE_mul_reg_2__15_ ( .D(PE_N47), .CK(clk), .Q(PE_mul[111]) );
  QDFFS PE_mul_reg_1__0_ ( .D(PE_N16), .CK(clk), .Q(PE_mul[112]) );
  QDFFS PE_mul_reg_1__1_ ( .D(PE_N17), .CK(clk), .Q(PE_mul[113]) );
  QDFFS PE_mul_reg_1__2_ ( .D(PE_N18), .CK(clk), .Q(PE_mul[114]) );
  QDFFS PE_mul_reg_1__3_ ( .D(PE_N19), .CK(clk), .Q(PE_mul[115]) );
  QDFFS PE_mul_reg_1__4_ ( .D(PE_N20), .CK(clk), .Q(PE_mul[116]) );
  QDFFS PE_mul_reg_1__5_ ( .D(PE_N21), .CK(clk), .Q(PE_mul[117]) );
  QDFFS PE_mul_reg_1__6_ ( .D(PE_N22), .CK(clk), .Q(PE_mul[118]) );
  QDFFS PE_mul_reg_1__7_ ( .D(PE_N23), .CK(clk), .Q(PE_mul[119]) );
  QDFFS PE_mul_reg_1__8_ ( .D(PE_N24), .CK(clk), .Q(PE_mul[120]) );
  QDFFS PE_mul_reg_1__9_ ( .D(PE_N25), .CK(clk), .Q(PE_mul[121]) );
  QDFFS PE_mul_reg_1__10_ ( .D(PE_N26), .CK(clk), .Q(PE_mul[122]) );
  QDFFS PE_mul_reg_1__11_ ( .D(PE_N27), .CK(clk), .Q(PE_mul[123]) );
  QDFFS PE_mul_reg_1__12_ ( .D(PE_N28), .CK(clk), .Q(PE_mul[124]) );
  QDFFS PE_mul_reg_1__13_ ( .D(PE_N29), .CK(clk), .Q(PE_mul[125]) );
  QDFFS PE_mul_reg_1__14_ ( .D(PE_N30), .CK(clk), .Q(PE_mul[126]) );
  QDFFS PE_mul_reg_1__15_ ( .D(PE_N31), .CK(clk), .Q(PE_mul[127]) );
  QDFFS PE_mul_reg_0__0_ ( .D(PE_N0), .CK(clk), .Q(PE_mul[128]) );
  QDFFS PE_mul_reg_0__1_ ( .D(PE_N1), .CK(clk), .Q(PE_mul[129]) );
  QDFFS PE_mul_reg_0__2_ ( .D(PE_N2), .CK(clk), .Q(PE_mul[130]) );
  QDFFS PE_mul_reg_0__3_ ( .D(PE_N3), .CK(clk), .Q(PE_mul[131]) );
  QDFFS PE_mul_reg_0__4_ ( .D(PE_N4), .CK(clk), .Q(PE_mul[132]) );
  QDFFS PE_mul_reg_0__5_ ( .D(PE_N5), .CK(clk), .Q(PE_mul[133]) );
  QDFFS PE_mul_reg_0__6_ ( .D(PE_N6), .CK(clk), .Q(PE_mul[134]) );
  QDFFS PE_mul_reg_0__7_ ( .D(PE_N7), .CK(clk), .Q(PE_mul[135]) );
  QDFFS PE_mul_reg_0__8_ ( .D(PE_N8), .CK(clk), .Q(PE_mul[136]) );
  QDFFS PE_mul_reg_0__9_ ( .D(PE_N9), .CK(clk), .Q(PE_mul[137]) );
  QDFFS PE_mul_reg_0__10_ ( .D(PE_N10), .CK(clk), .Q(PE_mul[138]) );
  QDFFS PE_mul_reg_0__11_ ( .D(PE_N11), .CK(clk), .Q(PE_mul[139]) );
  QDFFS PE_mul_reg_0__12_ ( .D(PE_N12), .CK(clk), .Q(PE_mul[140]) );
  QDFFS PE_mul_reg_0__13_ ( .D(PE_N13), .CK(clk), .Q(PE_mul[141]) );
  QDFFS PE_mul_reg_0__14_ ( .D(PE_N14), .CK(clk), .Q(PE_mul[142]) );
  QDFFS PE_mul_reg_0__15_ ( .D(PE_N15), .CK(clk), .Q(PE_mul[143]) );
  QDFFS m0_DO_reg_0_ ( .D(m0_DO_reg[0]), .CK(clk), .Q(gray_max_out[0]) );
  QDFFS m0_DO_reg_1_ ( .D(m0_DO_reg[1]), .CK(clk), .Q(gray_max_out[1]) );
  QDFFS m0_DO_reg_2_ ( .D(m0_DO_reg[2]), .CK(clk), .Q(gray_max_out[2]) );
  QDFFS m0_DO_reg_3_ ( .D(m0_DO_reg[3]), .CK(clk), .Q(gray_max_out[3]) );
  QDFFS m0_DO_reg_4_ ( .D(m0_DO_reg[4]), .CK(clk), .Q(gray_max_out[4]) );
  QDFFS m0_DO_reg_5_ ( .D(m0_DO_reg[5]), .CK(clk), .Q(gray_max_out[5]) );
  QDFFS m0_DO_reg_6_ ( .D(m0_DO_reg[6]), .CK(clk), .Q(gray_max_out[6]) );
  QDFFS m0_DO_reg_7_ ( .D(m0_DO_reg[7]), .CK(clk), .Q(gray_max_out[7]) );
  QDFFS m2_DO_reg_0_ ( .D(m2_DO_reg[0]), .CK(clk), .Q(gray_weight_out[0]) );
  QDFFS m2_DO_reg_1_ ( .D(m2_DO_reg[1]), .CK(clk), .Q(gray_weight_out[1]) );
  QDFFS m2_DO_reg_2_ ( .D(m2_DO_reg[2]), .CK(clk), .Q(gray_weight_out[2]) );
  QDFFS m2_DO_reg_3_ ( .D(m2_DO_reg[3]), .CK(clk), .Q(gray_weight_out[3]) );
  QDFFS m2_DO_reg_4_ ( .D(m2_DO_reg[4]), .CK(clk), .Q(gray_weight_out[4]) );
  QDFFS m2_DO_reg_5_ ( .D(m2_DO_reg[5]), .CK(clk), .Q(gray_weight_out[5]) );
  QDFFS m2_DO_reg_6_ ( .D(m2_DO_reg[6]), .CK(clk), .Q(gray_weight_out[6]) );
  QDFFS m2_DO_reg_7_ ( .D(m2_DO_reg[7]), .CK(clk), .Q(gray_weight_out[7]) );
  QDFFS m1_DO_reg_0_ ( .D(m1_DO_reg[0]), .CK(clk), .Q(gray_avg_out[0]) );
  QDFFS A67_shift_reg_0__0_ ( .D(n11261), .CK(clk), .Q(A67_shift[0]) );
  QDFFS A67_shift_reg_1__0_ ( .D(n11260), .CK(clk), .Q(A67_shift[8]) );
  QDFFS A67_shift_reg_2__0_ ( .D(n11259), .CK(clk), .Q(A67_shift[16]) );
  QDFFS A67_shift_reg_3__0_ ( .D(n11258), .CK(clk), .Q(A67_shift[24]) );
  QDFFS A67_shift_reg_4__0_ ( .D(n11257), .CK(clk), .Q(A67_shift[32]) );
  QDFFS A67_shift_reg_5__0_ ( .D(n11256), .CK(clk), .Q(A67_shift[40]) );
  QDFFS A67_shift_reg_6__0_ ( .D(n11255), .CK(clk), .Q(A67_shift[48]) );
  QDFFS A67_shift_reg_7__0_ ( .D(n11254), .CK(clk), .Q(A67_shift[56]) );
  QDFFS A67_shift_reg_8__0_ ( .D(n11253), .CK(clk), .Q(A67_shift[64]) );
  QDFFS A67_shift_reg_9__0_ ( .D(n11252), .CK(clk), .Q(A67_shift[72]) );
  QDFFS A67_shift_reg_10__0_ ( .D(n11251), .CK(clk), .Q(A67_shift[80]) );
  QDFFS A67_shift_reg_11__0_ ( .D(n11250), .CK(clk), .Q(A67_shift[88]) );
  QDFFS A67_shift_reg_12__0_ ( .D(n11249), .CK(clk), .Q(A67_shift[96]) );
  QDFFS A67_shift_reg_13__0_ ( .D(n11248), .CK(clk), .Q(A67_shift[104]) );
  QDFFS A67_shift_reg_14__0_ ( .D(n11247), .CK(clk), .Q(A67_shift[112]) );
  QDFFS A67_shift_reg_15__0_ ( .D(n11246), .CK(clk), .Q(A67_shift[120]) );
  QDFFS A67_shift_reg_16__0_ ( .D(n11245), .CK(clk), .Q(A67_shift[128]) );
  QDFFS A67_shift_reg_17__0_ ( .D(n11244), .CK(clk), .Q(A67_shift[136]) );
  QDFFS A67_shift_reg_18__0_ ( .D(n11243), .CK(clk), .Q(A67_shift[144]) );
  QDFFS A67_shift_reg_19__0_ ( .D(n11242), .CK(clk), .Q(A67_shift[152]) );
  QDFFS A67_shift_reg_20__0_ ( .D(n11241), .CK(clk), .Q(A67_shift[160]) );
  QDFFS A67_shift_reg_21__0_ ( .D(n11240), .CK(clk), .Q(A67_shift[168]) );
  QDFFS A67_shift_reg_22__0_ ( .D(n11239), .CK(clk), .Q(A67_shift[176]) );
  QDFFS A67_shift_reg_23__0_ ( .D(n11238), .CK(clk), .Q(A67_shift[184]) );
  QDFFS A67_shift_reg_24__0_ ( .D(n11237), .CK(clk), .Q(A67_shift[192]) );
  QDFFS A67_shift_reg_25__0_ ( .D(n11236), .CK(clk), .Q(A67_shift[200]) );
  QDFFS A67_shift_reg_26__0_ ( .D(n11235), .CK(clk), .Q(A67_shift[208]) );
  QDFFS A67_shift_reg_27__0_ ( .D(n11234), .CK(clk), .Q(A67_shift[216]) );
  QDFFS A67_shift_reg_28__0_ ( .D(n11233), .CK(clk), .Q(A67_shift[224]) );
  QDFFS A67_shift_reg_29__0_ ( .D(n11232), .CK(clk), .Q(A67_shift[232]) );
  QDFFS A67_shift_reg_30__0_ ( .D(n11231), .CK(clk), .Q(A67_shift[240]) );
  QDFFS A67_shift_reg_31__0_ ( .D(n11229), .CK(clk), .Q(A67_shift[248]) );
  QDFFS m1_DO_reg_1_ ( .D(m1_DO_reg[1]), .CK(clk), .Q(gray_avg_out[1]) );
  QDFFS A67_shift_reg_1__1_ ( .D(n11292), .CK(clk), .Q(A67_shift[9]) );
  QDFFS A67_shift_reg_2__1_ ( .D(n11291), .CK(clk), .Q(A67_shift[17]) );
  QDFFS A67_shift_reg_3__1_ ( .D(n11290), .CK(clk), .Q(A67_shift[25]) );
  QDFFS A67_shift_reg_4__1_ ( .D(n11289), .CK(clk), .Q(A67_shift[33]) );
  QDFFS A67_shift_reg_5__1_ ( .D(n11288), .CK(clk), .Q(A67_shift[41]) );
  QDFFS A67_shift_reg_6__1_ ( .D(n11287), .CK(clk), .Q(A67_shift[49]) );
  QDFFS A67_shift_reg_7__1_ ( .D(n11286), .CK(clk), .Q(A67_shift[57]) );
  QDFFS A67_shift_reg_8__1_ ( .D(n11285), .CK(clk), .Q(A67_shift[65]) );
  QDFFS A67_shift_reg_9__1_ ( .D(n11284), .CK(clk), .Q(A67_shift[73]) );
  QDFFS A67_shift_reg_10__1_ ( .D(n11283), .CK(clk), .Q(A67_shift[81]) );
  QDFFS A67_shift_reg_11__1_ ( .D(n11282), .CK(clk), .Q(A67_shift[89]) );
  QDFFS A67_shift_reg_12__1_ ( .D(n11281), .CK(clk), .Q(A67_shift[97]) );
  QDFFS A67_shift_reg_13__1_ ( .D(n11280), .CK(clk), .Q(A67_shift[105]) );
  QDFFS A67_shift_reg_14__1_ ( .D(n11279), .CK(clk), .Q(A67_shift[113]) );
  QDFFS A67_shift_reg_15__1_ ( .D(n11278), .CK(clk), .Q(A67_shift[121]) );
  QDFFS A67_shift_reg_16__1_ ( .D(n11277), .CK(clk), .Q(A67_shift[129]) );
  QDFFS A67_shift_reg_17__1_ ( .D(n11276), .CK(clk), .Q(A67_shift[137]) );
  QDFFS A67_shift_reg_18__1_ ( .D(n11275), .CK(clk), .Q(A67_shift[145]) );
  QDFFS A67_shift_reg_19__1_ ( .D(n11274), .CK(clk), .Q(A67_shift[153]) );
  QDFFS A67_shift_reg_20__1_ ( .D(n11273), .CK(clk), .Q(A67_shift[161]) );
  QDFFS A67_shift_reg_21__1_ ( .D(n11272), .CK(clk), .Q(A67_shift[169]) );
  QDFFS A67_shift_reg_22__1_ ( .D(n11271), .CK(clk), .Q(A67_shift[177]) );
  QDFFS A67_shift_reg_23__1_ ( .D(n11270), .CK(clk), .Q(A67_shift[185]) );
  QDFFS A67_shift_reg_24__1_ ( .D(n11269), .CK(clk), .Q(A67_shift[193]) );
  QDFFS A67_shift_reg_25__1_ ( .D(n11268), .CK(clk), .Q(A67_shift[201]) );
  QDFFS A67_shift_reg_26__1_ ( .D(n11267), .CK(clk), .Q(A67_shift[209]) );
  QDFFS A67_shift_reg_27__1_ ( .D(n11266), .CK(clk), .Q(A67_shift[217]) );
  QDFFS A67_shift_reg_28__1_ ( .D(n11265), .CK(clk), .Q(A67_shift[225]) );
  QDFFS A67_shift_reg_29__1_ ( .D(n11264), .CK(clk), .Q(A67_shift[233]) );
  QDFFS A67_shift_reg_30__1_ ( .D(n11263), .CK(clk), .Q(A67_shift[241]) );
  QDFFS A67_shift_reg_31__1_ ( .D(n11262), .CK(clk), .Q(A67_shift[249]) );
  QDFFS m1_DO_reg_2_ ( .D(m1_DO_reg[2]), .CK(clk), .Q(gray_avg_out[2]) );
  QDFFS A67_shift_reg_1__2_ ( .D(n11324), .CK(clk), .Q(A67_shift[10]) );
  QDFFS A67_shift_reg_2__2_ ( .D(n11323), .CK(clk), .Q(A67_shift[18]) );
  QDFFS A67_shift_reg_3__2_ ( .D(n11322), .CK(clk), .Q(A67_shift[26]) );
  QDFFS A67_shift_reg_4__2_ ( .D(n11321), .CK(clk), .Q(A67_shift[34]) );
  QDFFS A67_shift_reg_5__2_ ( .D(n11320), .CK(clk), .Q(A67_shift[42]) );
  QDFFS A67_shift_reg_6__2_ ( .D(n11319), .CK(clk), .Q(A67_shift[50]) );
  QDFFS A67_shift_reg_7__2_ ( .D(n11318), .CK(clk), .Q(A67_shift[58]) );
  QDFFS A67_shift_reg_8__2_ ( .D(n11317), .CK(clk), .Q(A67_shift[66]) );
  QDFFS A67_shift_reg_9__2_ ( .D(n11316), .CK(clk), .Q(A67_shift[74]) );
  QDFFS A67_shift_reg_10__2_ ( .D(n11315), .CK(clk), .Q(A67_shift[82]) );
  QDFFS A67_shift_reg_11__2_ ( .D(n11314), .CK(clk), .Q(A67_shift[90]) );
  QDFFS A67_shift_reg_12__2_ ( .D(n11313), .CK(clk), .Q(A67_shift[98]) );
  QDFFS A67_shift_reg_13__2_ ( .D(n11312), .CK(clk), .Q(A67_shift[106]) );
  QDFFS A67_shift_reg_14__2_ ( .D(n11311), .CK(clk), .Q(A67_shift[114]) );
  QDFFS A67_shift_reg_15__2_ ( .D(n11310), .CK(clk), .Q(A67_shift[122]) );
  QDFFS A67_shift_reg_16__2_ ( .D(n11309), .CK(clk), .Q(A67_shift[130]) );
  QDFFS A67_shift_reg_17__2_ ( .D(n11308), .CK(clk), .Q(A67_shift[138]) );
  QDFFS A67_shift_reg_18__2_ ( .D(n11307), .CK(clk), .Q(A67_shift[146]) );
  QDFFS A67_shift_reg_19__2_ ( .D(n11306), .CK(clk), .Q(A67_shift[154]) );
  QDFFS A67_shift_reg_20__2_ ( .D(n11305), .CK(clk), .Q(A67_shift[162]) );
  QDFFS A67_shift_reg_21__2_ ( .D(n11304), .CK(clk), .Q(A67_shift[170]) );
  QDFFS A67_shift_reg_22__2_ ( .D(n11303), .CK(clk), .Q(A67_shift[178]) );
  QDFFS A67_shift_reg_23__2_ ( .D(n11302), .CK(clk), .Q(A67_shift[186]) );
  QDFFS A67_shift_reg_24__2_ ( .D(n11301), .CK(clk), .Q(A67_shift[194]) );
  QDFFS A67_shift_reg_25__2_ ( .D(n11300), .CK(clk), .Q(A67_shift[202]) );
  QDFFS A67_shift_reg_26__2_ ( .D(n11299), .CK(clk), .Q(A67_shift[210]) );
  QDFFS A67_shift_reg_27__2_ ( .D(n11298), .CK(clk), .Q(A67_shift[218]) );
  QDFFS A67_shift_reg_28__2_ ( .D(n11297), .CK(clk), .Q(A67_shift[226]) );
  QDFFS A67_shift_reg_29__2_ ( .D(n11296), .CK(clk), .Q(A67_shift[234]) );
  QDFFS A67_shift_reg_30__2_ ( .D(n11295), .CK(clk), .Q(A67_shift[242]) );
  QDFFS A67_shift_reg_31__2_ ( .D(n11294), .CK(clk), .Q(A67_shift[250]) );
  QDFFS m1_DO_reg_3_ ( .D(m1_DO_reg[3]), .CK(clk), .Q(gray_avg_out[3]) );
  QDFFS A67_shift_reg_1__3_ ( .D(n11356), .CK(clk), .Q(A67_shift[11]) );
  QDFFS A67_shift_reg_2__3_ ( .D(n11355), .CK(clk), .Q(A67_shift[19]) );
  QDFFS A67_shift_reg_3__3_ ( .D(n11354), .CK(clk), .Q(A67_shift[27]) );
  QDFFS A67_shift_reg_4__3_ ( .D(n11353), .CK(clk), .Q(A67_shift[35]) );
  QDFFS A67_shift_reg_5__3_ ( .D(n11352), .CK(clk), .Q(A67_shift[43]) );
  QDFFS A67_shift_reg_6__3_ ( .D(n11351), .CK(clk), .Q(A67_shift[51]) );
  QDFFS A67_shift_reg_7__3_ ( .D(n11350), .CK(clk), .Q(A67_shift[59]) );
  QDFFS A67_shift_reg_8__3_ ( .D(n11349), .CK(clk), .Q(A67_shift[67]) );
  QDFFS A67_shift_reg_9__3_ ( .D(n11348), .CK(clk), .Q(A67_shift[75]) );
  QDFFS A67_shift_reg_10__3_ ( .D(n11347), .CK(clk), .Q(A67_shift[83]) );
  QDFFS A67_shift_reg_11__3_ ( .D(n11346), .CK(clk), .Q(A67_shift[91]) );
  QDFFS A67_shift_reg_12__3_ ( .D(n11345), .CK(clk), .Q(A67_shift[99]) );
  QDFFS A67_shift_reg_13__3_ ( .D(n11344), .CK(clk), .Q(A67_shift[107]) );
  QDFFS A67_shift_reg_14__3_ ( .D(n11343), .CK(clk), .Q(A67_shift[115]) );
  QDFFS A67_shift_reg_15__3_ ( .D(n11342), .CK(clk), .Q(A67_shift[123]) );
  QDFFS A67_shift_reg_16__3_ ( .D(n11341), .CK(clk), .Q(A67_shift[131]) );
  QDFFS A67_shift_reg_17__3_ ( .D(n11340), .CK(clk), .Q(A67_shift[139]) );
  QDFFS A67_shift_reg_18__3_ ( .D(n11339), .CK(clk), .Q(A67_shift[147]) );
  QDFFS A67_shift_reg_19__3_ ( .D(n11338), .CK(clk), .Q(A67_shift[155]) );
  QDFFS A67_shift_reg_20__3_ ( .D(n11337), .CK(clk), .Q(A67_shift[163]) );
  QDFFS A67_shift_reg_21__3_ ( .D(n11336), .CK(clk), .Q(A67_shift[171]) );
  QDFFS A67_shift_reg_22__3_ ( .D(n11335), .CK(clk), .Q(A67_shift[179]) );
  QDFFS A67_shift_reg_23__3_ ( .D(n11334), .CK(clk), .Q(A67_shift[187]) );
  QDFFS A67_shift_reg_24__3_ ( .D(n11333), .CK(clk), .Q(A67_shift[195]) );
  QDFFS A67_shift_reg_25__3_ ( .D(n11332), .CK(clk), .Q(A67_shift[203]) );
  QDFFS A67_shift_reg_26__3_ ( .D(n11331), .CK(clk), .Q(A67_shift[211]) );
  QDFFS A67_shift_reg_27__3_ ( .D(n11330), .CK(clk), .Q(A67_shift[219]) );
  QDFFS A67_shift_reg_28__3_ ( .D(n11329), .CK(clk), .Q(A67_shift[227]) );
  QDFFS A67_shift_reg_29__3_ ( .D(n11328), .CK(clk), .Q(A67_shift[235]) );
  QDFFS A67_shift_reg_30__3_ ( .D(n11327), .CK(clk), .Q(A67_shift[243]) );
  QDFFS A67_shift_reg_31__3_ ( .D(n11326), .CK(clk), .Q(A67_shift[251]) );
  QDFFS m1_DO_reg_4_ ( .D(m1_DO_reg[4]), .CK(clk), .Q(gray_avg_out[4]) );
  QDFFS A67_shift_reg_0__4_ ( .D(n11389), .CK(clk), .Q(A67_shift[4]) );
  QDFFS A67_shift_reg_1__4_ ( .D(n11388), .CK(clk), .Q(A67_shift[12]) );
  QDFFS A67_shift_reg_2__4_ ( .D(n11387), .CK(clk), .Q(A67_shift[20]) );
  QDFFS A67_shift_reg_3__4_ ( .D(n11386), .CK(clk), .Q(A67_shift[28]) );
  QDFFS A67_shift_reg_4__4_ ( .D(n11385), .CK(clk), .Q(A67_shift[36]) );
  QDFFS A67_shift_reg_5__4_ ( .D(n11384), .CK(clk), .Q(A67_shift[44]) );
  QDFFS A67_shift_reg_6__4_ ( .D(n11383), .CK(clk), .Q(A67_shift[52]) );
  QDFFS A67_shift_reg_7__4_ ( .D(n11382), .CK(clk), .Q(A67_shift[60]) );
  QDFFS A67_shift_reg_8__4_ ( .D(n11381), .CK(clk), .Q(A67_shift[68]) );
  QDFFS A67_shift_reg_9__4_ ( .D(n11380), .CK(clk), .Q(A67_shift[76]) );
  QDFFS A67_shift_reg_10__4_ ( .D(n11379), .CK(clk), .Q(A67_shift[84]) );
  QDFFS A67_shift_reg_11__4_ ( .D(n11378), .CK(clk), .Q(A67_shift[92]) );
  QDFFS A67_shift_reg_12__4_ ( .D(n11377), .CK(clk), .Q(A67_shift[100]) );
  QDFFS A67_shift_reg_13__4_ ( .D(n11376), .CK(clk), .Q(A67_shift[108]) );
  QDFFS A67_shift_reg_14__4_ ( .D(n11375), .CK(clk), .Q(A67_shift[116]) );
  QDFFS A67_shift_reg_15__4_ ( .D(n11374), .CK(clk), .Q(A67_shift[124]) );
  QDFFS A67_shift_reg_16__4_ ( .D(n11373), .CK(clk), .Q(A67_shift[132]) );
  QDFFS A67_shift_reg_17__4_ ( .D(n11372), .CK(clk), .Q(A67_shift[140]) );
  QDFFS A67_shift_reg_18__4_ ( .D(n11371), .CK(clk), .Q(A67_shift[148]) );
  QDFFS A67_shift_reg_19__4_ ( .D(n11370), .CK(clk), .Q(A67_shift[156]) );
  QDFFS A67_shift_reg_20__4_ ( .D(n11369), .CK(clk), .Q(A67_shift[164]) );
  QDFFS A67_shift_reg_21__4_ ( .D(n11368), .CK(clk), .Q(A67_shift[172]) );
  QDFFS A67_shift_reg_22__4_ ( .D(n11367), .CK(clk), .Q(A67_shift[180]) );
  QDFFS A67_shift_reg_23__4_ ( .D(n11366), .CK(clk), .Q(A67_shift[188]) );
  QDFFS A67_shift_reg_24__4_ ( .D(n11365), .CK(clk), .Q(A67_shift[196]) );
  QDFFS A67_shift_reg_25__4_ ( .D(n11364), .CK(clk), .Q(A67_shift[204]) );
  QDFFS A67_shift_reg_26__4_ ( .D(n11363), .CK(clk), .Q(A67_shift[212]) );
  QDFFS A67_shift_reg_27__4_ ( .D(n11362), .CK(clk), .Q(A67_shift[220]) );
  QDFFS A67_shift_reg_28__4_ ( .D(n11361), .CK(clk), .Q(A67_shift[228]) );
  QDFFS A67_shift_reg_29__4_ ( .D(n11360), .CK(clk), .Q(A67_shift[236]) );
  QDFFS A67_shift_reg_30__4_ ( .D(n11359), .CK(clk), .Q(A67_shift[244]) );
  QDFFS A67_shift_reg_31__4_ ( .D(n11358), .CK(clk), .Q(A67_shift[252]) );
  QDFFS m1_DO_reg_5_ ( .D(m1_DO_reg[5]), .CK(clk), .Q(gray_avg_out[5]) );
  QDFFS A67_shift_reg_1__5_ ( .D(n11420), .CK(clk), .Q(A67_shift[13]) );
  QDFFS A67_shift_reg_2__5_ ( .D(n11419), .CK(clk), .Q(A67_shift[21]) );
  QDFFS A67_shift_reg_3__5_ ( .D(n11418), .CK(clk), .Q(A67_shift[29]) );
  QDFFS A67_shift_reg_4__5_ ( .D(n11417), .CK(clk), .Q(A67_shift[37]) );
  QDFFS A67_shift_reg_5__5_ ( .D(n11416), .CK(clk), .Q(A67_shift[45]) );
  QDFFS A67_shift_reg_6__5_ ( .D(n11415), .CK(clk), .Q(A67_shift[53]) );
  QDFFS A67_shift_reg_7__5_ ( .D(n11414), .CK(clk), .Q(A67_shift[61]) );
  QDFFS A67_shift_reg_8__5_ ( .D(n11413), .CK(clk), .Q(A67_shift[69]) );
  QDFFS A67_shift_reg_9__5_ ( .D(n11412), .CK(clk), .Q(A67_shift[77]) );
  QDFFS A67_shift_reg_10__5_ ( .D(n11411), .CK(clk), .Q(A67_shift[85]) );
  QDFFS A67_shift_reg_11__5_ ( .D(n11410), .CK(clk), .Q(A67_shift[93]) );
  QDFFS A67_shift_reg_12__5_ ( .D(n11409), .CK(clk), .Q(A67_shift[101]) );
  QDFFS A67_shift_reg_13__5_ ( .D(n11408), .CK(clk), .Q(A67_shift[109]) );
  QDFFS A67_shift_reg_14__5_ ( .D(n11407), .CK(clk), .Q(A67_shift[117]) );
  QDFFS A67_shift_reg_15__5_ ( .D(n11406), .CK(clk), .Q(A67_shift[125]) );
  QDFFS A67_shift_reg_16__5_ ( .D(n11405), .CK(clk), .Q(A67_shift[133]) );
  QDFFS A67_shift_reg_17__5_ ( .D(n11404), .CK(clk), .Q(A67_shift[141]) );
  QDFFS A67_shift_reg_18__5_ ( .D(n11403), .CK(clk), .Q(A67_shift[149]) );
  QDFFS A67_shift_reg_19__5_ ( .D(n11402), .CK(clk), .Q(A67_shift[157]) );
  QDFFS A67_shift_reg_20__5_ ( .D(n11401), .CK(clk), .Q(A67_shift[165]) );
  QDFFS A67_shift_reg_21__5_ ( .D(n11400), .CK(clk), .Q(A67_shift[173]) );
  QDFFS A67_shift_reg_22__5_ ( .D(n11399), .CK(clk), .Q(A67_shift[181]) );
  QDFFS A67_shift_reg_23__5_ ( .D(n11398), .CK(clk), .Q(A67_shift[189]) );
  QDFFS A67_shift_reg_24__5_ ( .D(n11397), .CK(clk), .Q(A67_shift[197]) );
  QDFFS A67_shift_reg_25__5_ ( .D(n11396), .CK(clk), .Q(A67_shift[205]) );
  QDFFS A67_shift_reg_26__5_ ( .D(n11395), .CK(clk), .Q(A67_shift[213]) );
  QDFFS A67_shift_reg_27__5_ ( .D(n11394), .CK(clk), .Q(A67_shift[221]) );
  QDFFS A67_shift_reg_28__5_ ( .D(n11393), .CK(clk), .Q(A67_shift[229]) );
  QDFFS A67_shift_reg_29__5_ ( .D(n11392), .CK(clk), .Q(A67_shift[237]) );
  QDFFS A67_shift_reg_30__5_ ( .D(n11391), .CK(clk), .Q(A67_shift[245]) );
  QDFFS A67_shift_reg_31__5_ ( .D(n11390), .CK(clk), .Q(A67_shift[253]) );
  QDFFS m1_DO_reg_6_ ( .D(m1_DO_reg[6]), .CK(clk), .Q(gray_avg_out[6]) );
  QDFFS A67_shift_reg_1__6_ ( .D(n11452), .CK(clk), .Q(A67_shift[14]) );
  QDFFS A67_shift_reg_2__6_ ( .D(n11451), .CK(clk), .Q(A67_shift[22]) );
  QDFFS A67_shift_reg_3__6_ ( .D(n11450), .CK(clk), .Q(A67_shift[30]) );
  QDFFS A67_shift_reg_4__6_ ( .D(n11449), .CK(clk), .Q(A67_shift[38]) );
  QDFFS A67_shift_reg_5__6_ ( .D(n11448), .CK(clk), .Q(A67_shift[46]) );
  QDFFS A67_shift_reg_6__6_ ( .D(n11447), .CK(clk), .Q(A67_shift[54]) );
  QDFFS A67_shift_reg_7__6_ ( .D(n11446), .CK(clk), .Q(A67_shift[62]) );
  QDFFS A67_shift_reg_8__6_ ( .D(n11445), .CK(clk), .Q(A67_shift[70]) );
  QDFFS A67_shift_reg_9__6_ ( .D(n11444), .CK(clk), .Q(A67_shift[78]) );
  QDFFS A67_shift_reg_10__6_ ( .D(n11443), .CK(clk), .Q(A67_shift[86]) );
  QDFFS A67_shift_reg_11__6_ ( .D(n11442), .CK(clk), .Q(A67_shift[94]) );
  QDFFS A67_shift_reg_12__6_ ( .D(n11441), .CK(clk), .Q(A67_shift[102]) );
  QDFFS A67_shift_reg_13__6_ ( .D(n11440), .CK(clk), .Q(A67_shift[110]) );
  QDFFS A67_shift_reg_14__6_ ( .D(n11439), .CK(clk), .Q(A67_shift[118]) );
  QDFFS A67_shift_reg_15__6_ ( .D(n11438), .CK(clk), .Q(A67_shift[126]) );
  QDFFS A67_shift_reg_16__6_ ( .D(n11437), .CK(clk), .Q(A67_shift[134]) );
  QDFFS A67_shift_reg_17__6_ ( .D(n11436), .CK(clk), .Q(A67_shift[142]) );
  QDFFS A67_shift_reg_18__6_ ( .D(n11435), .CK(clk), .Q(A67_shift[150]) );
  QDFFS A67_shift_reg_19__6_ ( .D(n11434), .CK(clk), .Q(A67_shift[158]) );
  QDFFS A67_shift_reg_20__6_ ( .D(n11433), .CK(clk), .Q(A67_shift[166]) );
  QDFFS A67_shift_reg_21__6_ ( .D(n11432), .CK(clk), .Q(A67_shift[174]) );
  QDFFS A67_shift_reg_22__6_ ( .D(n11431), .CK(clk), .Q(A67_shift[182]) );
  QDFFS A67_shift_reg_23__6_ ( .D(n11430), .CK(clk), .Q(A67_shift[190]) );
  QDFFS A67_shift_reg_24__6_ ( .D(n11429), .CK(clk), .Q(A67_shift[198]) );
  QDFFS A67_shift_reg_25__6_ ( .D(n11428), .CK(clk), .Q(A67_shift[206]) );
  QDFFS A67_shift_reg_26__6_ ( .D(n11427), .CK(clk), .Q(A67_shift[214]) );
  QDFFS A67_shift_reg_27__6_ ( .D(n11426), .CK(clk), .Q(A67_shift[222]) );
  QDFFS A67_shift_reg_28__6_ ( .D(n11425), .CK(clk), .Q(A67_shift[230]) );
  QDFFS A67_shift_reg_29__6_ ( .D(n11424), .CK(clk), .Q(A67_shift[238]) );
  QDFFS A67_shift_reg_30__6_ ( .D(n11423), .CK(clk), .Q(A67_shift[246]) );
  QDFFS A67_shift_reg_31__6_ ( .D(n11422), .CK(clk), .Q(A67_shift[254]) );
  QDFFS m1_DO_reg_7_ ( .D(m1_DO_reg[7]), .CK(clk), .Q(gray_avg_out[7]) );
  QDFFS A67_shift_reg_0__7_ ( .D(n11485), .CK(clk), .Q(A67_shift[7]) );
  QDFFS A67_shift_reg_1__7_ ( .D(n11484), .CK(clk), .Q(A67_shift[15]) );
  QDFFS A67_shift_reg_2__7_ ( .D(n11483), .CK(clk), .Q(A67_shift[23]) );
  QDFFS A67_shift_reg_3__7_ ( .D(n11482), .CK(clk), .Q(A67_shift[31]) );
  QDFFS A67_shift_reg_4__7_ ( .D(n11481), .CK(clk), .Q(A67_shift[39]) );
  QDFFS A67_shift_reg_5__7_ ( .D(n11480), .CK(clk), .Q(A67_shift[47]) );
  QDFFS A67_shift_reg_6__7_ ( .D(n11479), .CK(clk), .Q(A67_shift[55]) );
  QDFFS A67_shift_reg_7__7_ ( .D(n11478), .CK(clk), .Q(A67_shift[63]) );
  QDFFS A67_shift_reg_8__7_ ( .D(n11477), .CK(clk), .Q(A67_shift[71]) );
  QDFFS A67_shift_reg_9__7_ ( .D(n11476), .CK(clk), .Q(A67_shift[79]) );
  QDFFS A67_shift_reg_10__7_ ( .D(n11475), .CK(clk), .Q(A67_shift[87]) );
  QDFFS A67_shift_reg_11__7_ ( .D(n11474), .CK(clk), .Q(A67_shift[95]) );
  QDFFS A67_shift_reg_12__7_ ( .D(n11473), .CK(clk), .Q(A67_shift[103]) );
  QDFFS A67_shift_reg_13__7_ ( .D(n11472), .CK(clk), .Q(A67_shift[111]) );
  QDFFS A67_shift_reg_14__7_ ( .D(n11471), .CK(clk), .Q(A67_shift[119]) );
  QDFFS A67_shift_reg_15__7_ ( .D(n11470), .CK(clk), .Q(A67_shift[127]) );
  QDFFS A67_shift_reg_16__7_ ( .D(n11469), .CK(clk), .Q(A67_shift[135]) );
  QDFFS A67_shift_reg_17__7_ ( .D(n11468), .CK(clk), .Q(A67_shift[143]) );
  QDFFS A67_shift_reg_18__7_ ( .D(n11467), .CK(clk), .Q(A67_shift[151]) );
  QDFFS A67_shift_reg_19__7_ ( .D(n11466), .CK(clk), .Q(A67_shift[159]) );
  QDFFS A67_shift_reg_20__7_ ( .D(n11465), .CK(clk), .Q(A67_shift[167]) );
  QDFFS A67_shift_reg_21__7_ ( .D(n11464), .CK(clk), .Q(A67_shift[175]) );
  QDFFS A67_shift_reg_22__7_ ( .D(n11463), .CK(clk), .Q(A67_shift[183]) );
  QDFFS A67_shift_reg_23__7_ ( .D(n11462), .CK(clk), .Q(A67_shift[191]) );
  QDFFS A67_shift_reg_24__7_ ( .D(n11461), .CK(clk), .Q(A67_shift[199]) );
  QDFFS A67_shift_reg_25__7_ ( .D(n11460), .CK(clk), .Q(A67_shift[207]) );
  QDFFS A67_shift_reg_26__7_ ( .D(n11459), .CK(clk), .Q(A67_shift[215]) );
  QDFFS A67_shift_reg_27__7_ ( .D(n11458), .CK(clk), .Q(A67_shift[223]) );
  QDFFS A67_shift_reg_28__7_ ( .D(n11457), .CK(clk), .Q(A67_shift[231]) );
  QDFFS A67_shift_reg_29__7_ ( .D(n11456), .CK(clk), .Q(A67_shift[239]) );
  QDFFS A67_shift_reg_30__7_ ( .D(n11455), .CK(clk), .Q(A67_shift[247]) );
  QDFFS A67_shift_reg_31__7_ ( .D(n11454), .CK(clk), .Q(A67_shift[255]) );
  DFFSBN out_cnt_reg_1_ ( .D(n13683), .CK(clk), .SB(n30035), .Q(out_cnt[1]), 
        .QB(n30032) );
  DFFSBN out_cnt_reg_4_ ( .D(n13682), .CK(clk), .SB(n30035), .Q(out_cnt[4]), 
        .QB(n30033) );
  FA1S intadd_8_U8 ( .A(rgb_value[9]), .B(rgb_value[2]), .CI(rgb_value[18]), 
        .CO(intadd_8_n7), .S(gray_weight[0]) );
  FA1S intadd_8_U7 ( .A(intadd_8_B_1_), .B(rgb_value[3]), .CI(intadd_8_n7), 
        .CO(intadd_8_n6), .S(gray_weight[1]) );
  FA1S intadd_8_U6 ( .A(intadd_8_B_2_), .B(intadd_8_A_2_), .CI(intadd_8_n6), 
        .CO(intadd_8_n5), .S(gray_weight[2]) );
  FA1S intadd_8_U5 ( .A(intadd_8_B_3_), .B(intadd_8_A_3_), .CI(intadd_8_n5), 
        .CO(intadd_8_n4), .S(gray_weight[3]) );
  FA1S intadd_8_U4 ( .A(intadd_8_B_4_), .B(intadd_8_A_4_), .CI(intadd_8_n4), 
        .CO(intadd_8_n3), .S(gray_weight[4]) );
  FA1S intadd_8_U3 ( .A(intadd_8_B_5_), .B(intadd_8_A_5_), .CI(intadd_8_n3), 
        .CO(intadd_8_n2), .S(gray_weight[5]) );
  QDFFRBS c_s_reg_0_ ( .D(n30028), .CK(clk), .RB(n13805), .Q(c_s[0]) );
  QDFFRBS img_size_reg_2_ ( .D(n13642), .CK(clk), .RB(n13805), .Q(img_size[2])
         );
  QDFFRBS addr_reg_3_ ( .D(n13629), .CK(clk), .RB(n13805), .Q(addr[3]) );
  QDFFRBS addr_reg_6_ ( .D(n13626), .CK(clk), .RB(n13805), .Q(addr[6]) );
  QDFFRBS temp_cnt_reg_1_ ( .D(n13624), .CK(clk), .RB(n13805), .Q(temp_cnt[1])
         );
  QDFFRBT i_row_reg_1_ ( .D(n13608), .CK(clk), .RB(n13805), .Q(i_row[1]) );
  QDFFRBT i_row_reg_3_ ( .D(n13606), .CK(clk), .RB(n13805), .Q(i_row[3]) );
  QDFFRBS col_reg_1_ ( .D(n13621), .CK(clk), .RB(n13805), .Q(col[1]) );
  QDFFRBP i_col_reg_3_ ( .D(n13612), .CK(clk), .RB(n30034), .Q(i_col[3]) );
  QDFFRBN img_size_reg_0_ ( .D(n13689), .CK(clk), .RB(n13805), .Q(img_size[0])
         );
  QDFFRBT i_col_reg_1_ ( .D(n13610), .CK(clk), .RB(n30034), .Q(i_col[1]) );
  QDFFRBT img_size_reg_1_ ( .D(n13643), .CK(clk), .RB(n30034), .Q(img_size[1])
         );
  QDFFRBP i_col_reg_2_ ( .D(n13611), .CK(clk), .RB(n30034), .Q(i_col[2]) );
  QDFFP PE_mul_reg_4__15_ ( .D(PE_N79), .CK(clk), .Q(PE_mul[79]) );
  QDFFP PE_mul_reg_5__15_ ( .D(PE_N95), .CK(clk), .Q(PE_mul[63]) );
  QDFFP A67_shift_reg_0__2_ ( .D(n11325), .CK(clk), .Q(A67_shift[2]) );
  QDFFS A67_shift_reg_0__1_ ( .D(n11293), .CK(clk), .Q(A67_shift[1]) );
  QDFFS A67_shift_reg_0__5_ ( .D(n11421), .CK(clk), .Q(A67_shift[5]) );
  QDFFS A67_shift_reg_0__6_ ( .D(n11453), .CK(clk), .Q(A67_shift[6]) );
  QDFFP PE_mul_reg_3__15_ ( .D(PE_N63), .CK(clk), .Q(PE_mul[95]) );
  QDFFRBT i_row_reg_2_ ( .D(n13607), .CK(clk), .RB(n13805), .Q(i_row[2]) );
  QDFFS A67_shift_reg_0__3_ ( .D(n11357), .CK(clk), .Q(A67_shift[3]) );
  QDFFP img_reg_9__4__4_ ( .D(n12672), .CK(clk), .Q(img[860]) );
  QDFFP img_reg_9__1__5_ ( .D(n12649), .CK(clk), .Q(img[885]) );
  QDFFP img_reg_9__8__4_ ( .D(n12704), .CK(clk), .Q(img[828]) );
  QDFFP img_reg_5__7__5_ ( .D(n12185), .CK(clk), .Q(img[1349]) );
  QDFFP img_reg_3__7__5_ ( .D(n11929), .CK(clk), .Q(img[1605]) );
  QDFFP img_reg_4__3__5_ ( .D(n12023), .CK(clk), .Q(img[1509]) );
  QDFFP img_reg_3__3__5_ ( .D(n11896), .CK(clk), .Q(img[1637]) );
  QDFFP img_reg_7__6__5_ ( .D(n12431), .CK(clk), .Q(img[1101]) );
  QDFFP img_reg_6__6__5_ ( .D(n12305), .CK(clk), .Q(img[1229]) );
  QDFFP img_reg_4__5__3_ ( .D(n12041), .CK(clk), .Q(img[1491]) );
  QDFFRBT i_row_reg_0_ ( .D(n13609), .CK(clk), .RB(n13805), .Q(i_row[0]) );
  JKFRBN out_cnt_reg_0_ ( .J(n31997), .K(n31996), .CK(clk), .RB(n30035), .Q(
        n30030), .QB(out_cnt[0]) );
  JKFRBN act_ptr_reg_0_ ( .J(n30039), .K(n30036), .CK(clk), .RB(n30035), .Q(
        n30031), .QB(act_ptr[0]) );
  DFFN img_reg_4__7__5_ ( .D(n12055), .CK(clk), .Q(img[1477]), .QB(n30911) );
  DFFN img_reg_2__0__5_ ( .D(n11745), .CK(clk), .Q(img[1789]), .QB(n30809) );
  DFFN img_reg_3__5__3_ ( .D(n11911), .CK(clk), .Q(img[1619]), .QB(n31302) );
  DFFN img_reg_2__2__3_ ( .D(n11759), .CK(clk), .Q(img[1771]), .QB(n31295) );
  DFFN img_reg_2__6__0_ ( .D(n11796), .CK(clk), .Q(img[1736]), .QB(n31609) );
  DFFN img_reg_7__1__2_ ( .D(n12390), .CK(clk), .Q(img[1138]), .QB(n30581) );
  DFFN img_reg_0__2__2_ ( .D(n11502), .CK(clk), .Q(img[2026]), .QB(n30586) );
  DFFN img_reg_4__7__0_ ( .D(n12060), .CK(clk), .Q(img[1472]), .QB(n31514) );
  DFFN img_reg_3__6__6_ ( .D(n11918), .CK(clk), .Q(img[1614]), .QB(n30392) );
  DFFN img_reg_2__2__1_ ( .D(n11757), .CK(clk), .Q(img[1769]), .QB(n31159) );
  DFFN img_reg_4__6__4_ ( .D(n12048), .CK(clk), .Q(img[1484]), .QB(n31765) );
  DFFN img_reg_0__7__4_ ( .D(n11544), .CK(clk), .Q(img[1988]), .QB(n31865) );
  DFFN img_reg_14__5__5_ ( .D(n13319), .CK(clk), .Q(img[213]), .QB(n30928) );
  DFFN img_reg_14__10__5_ ( .D(n13361), .CK(clk), .Q(img[173]), .QB(n30927) );
  DFFN img_reg_7__14__5_ ( .D(n12495), .CK(clk), .Q(img[1037]), .QB(n30939) );
  DFFN img_reg_1__3__1_ ( .D(n11637), .CK(clk), .Q(img[1889]), .QB(n31041) );
  DFFN img_reg_12__10__5_ ( .D(n13105), .CK(clk), .Q(img[429]), .QB(n30931) );
  DFFN img_reg_12__5__5_ ( .D(n13063), .CK(clk), .Q(img[469]), .QB(n30932) );
  DFFN img_reg_4__7__6_ ( .D(n12054), .CK(clk), .Q(img[1478]), .QB(n30305) );
  DFFN img_reg_6__5__6_ ( .D(n12294), .CK(clk), .Q(img[1238]), .QB(n30500) );
  DFFN img_reg_0__6__6_ ( .D(n11538), .CK(clk), .Q(img[1998]), .QB(n30404) );
  DFFN img_reg_5__4__6_ ( .D(n12158), .CK(clk), .Q(img[1374]), .QB(n30416) );
  DFFN img_reg_6__3__6_ ( .D(n12278), .CK(clk), .Q(img[1254]), .QB(n30413) );
  DFFN img_reg_7__0__1_ ( .D(n12387), .CK(clk), .Q(img[1145]), .QB(n31064) );
  DFFN img_reg_2__7__1_ ( .D(n11803), .CK(clk), .Q(img[1729]), .QB(n31051) );
  DFFN img_reg_0__6__1_ ( .D(n11533), .CK(clk), .Q(img[1993]), .QB(n31175) );
  DFFN img_reg_5__2__1_ ( .D(n12147), .CK(clk), .Q(img[1385]), .QB(n31128) );
  DFFN img_reg_6__2__1_ ( .D(n12269), .CK(clk), .Q(img[1257]), .QB(n31124) );
  DFFN img_reg_3__5__7_ ( .D(n11915), .CK(clk), .Q(img[1623]), .QB(n30082) );
  DFFN img_reg_1__6__7_ ( .D(n11661), .CK(clk), .Q(img[1871]), .QB(n30072) );
  DFFN img_reg_7__4__7_ ( .D(n12413), .CK(clk), .Q(img[1119]), .QB(n30153) );
  DFFN img_reg_5__4__7_ ( .D(n12157), .CK(clk), .Q(img[1375]), .QB(n30110) );
  DFFN img_reg_1__0__6_ ( .D(n11614), .CK(clk), .Q(img[1918]), .QB(n30313) );
  DFFN img_reg_1__3__6_ ( .D(n11642), .CK(clk), .Q(img[1894]), .QB(n30311) );
  DFFN img_reg_1__1__6_ ( .D(n11626), .CK(clk), .Q(img[1910]), .QB(n30378) );
  DFFN img_reg_0__1__6_ ( .D(n11494), .CK(clk), .Q(img[2038]), .QB(n30406) );
  DFFN img_reg_2__3__1_ ( .D(n11771), .CK(clk), .Q(img[1761]), .QB(n31049) );
  DFFN img_reg_3__0__1_ ( .D(n11875), .CK(clk), .Q(img[1657]), .QB(n31060) );
  DFFN img_reg_2__2__7_ ( .D(n11763), .CK(clk), .Q(img[1775]), .QB(n30076) );
  DFFN img_reg_3__3__7_ ( .D(n11898), .CK(clk), .Q(img[1639]), .QB(n30150) );
  DFFN img_reg_2__1__7_ ( .D(n11749), .CK(clk), .Q(img[1783]), .QB(n30078) );
  DFFN img_reg_1__1__7_ ( .D(n11627), .CK(clk), .Q(img[1911]), .QB(n30070) );
  DFFN img_reg_0__1__7_ ( .D(n11493), .CK(clk), .Q(img[2039]), .QB(n30098) );
  DFFN img_reg_3__1__7_ ( .D(n11883), .CK(clk), .Q(img[1655]), .QB(n30086) );
  DFFN img_reg_12__1__0_ ( .D(n13036), .CK(clk), .Q(img[496]), .QB(n31654) );
  DFFN img_reg_14__1__0_ ( .D(n13292), .CK(clk), .Q(img[240]), .QB(n31650) );
  DFFN img_reg_3__6__4_ ( .D(n11920), .CK(clk), .Q(img[1612]), .QB(n31792) );
  DFFN img_reg_7__1__4_ ( .D(n12392), .CK(clk), .Q(img[1140]), .QB(n31794) );
  DFFN img_reg_2__7__4_ ( .D(n11800), .CK(clk), .Q(img[1732]), .QB(n31845) );
  DFFN img_reg_0__5__4_ ( .D(n11528), .CK(clk), .Q(img[2004]), .QB(n31798) );
  DFFN img_reg_7__3__4_ ( .D(n12408), .CK(clk), .Q(img[1124]), .QB(n31918) );
  DFFN img_reg_3__7__4_ ( .D(n11928), .CK(clk), .Q(img[1604]), .QB(n31853) );
  DFFN img_reg_0__2__4_ ( .D(n11504), .CK(clk), .Q(img[2028]), .QB(n31800) );
  DFFN img_reg_3__3__4_ ( .D(n11895), .CK(clk), .Q(img[1636]), .QB(n31850) );
  DFFN img_reg_2__3__4_ ( .D(n11768), .CK(clk), .Q(img[1764]), .QB(n31842) );
  DFFN img_reg_3__2__4_ ( .D(n11888), .CK(clk), .Q(img[1644]), .QB(n31788) );
  DFFN img_reg_12__1__3_ ( .D(n13033), .CK(clk), .Q(img[499]), .QB(n31407) );
  DFFN img_reg_14__1__3_ ( .D(n13289), .CK(clk), .Q(img[243]), .QB(n31403) );
  DFFN img_reg_0__14__1_ ( .D(n11597), .CK(clk), .Q(img[1929]), .QB(n31176) );
  DFFN img_reg_12__2__7_ ( .D(n13043), .CK(clk), .Q(img[495]), .QB(n30212) );
  DFFN img_reg_14__13__7_ ( .D(n13381), .CK(clk), .Q(img[151]), .QB(n30209) );
  DFFN img_reg_7__10__1_ ( .D(n12467), .CK(clk), .Q(img[1065]), .QB(n31172) );
  DFFN img_reg_3__13__1_ ( .D(n11973), .CK(clk), .Q(img[1553]), .QB(n31166) );
  DFFN img_reg_0__13__1_ ( .D(n11595), .CK(clk), .Q(img[1937]), .QB(n31178) );
  DFFN img_reg_2__6__5_ ( .D(n11793), .CK(clk), .Q(img[1741]), .QB(n30868) );
  DFFN img_reg_4__6__5_ ( .D(n12049), .CK(clk), .Q(img[1485]), .QB(n30964) );
  DFFN img_reg_0__7__5_ ( .D(n11543), .CK(clk), .Q(img[1989]), .QB(n30825) );
  DFFN img_reg_6__5__5_ ( .D(n12295), .CK(clk), .Q(img[1237]), .QB(n30837) );
  DFFN img_reg_7__5__5_ ( .D(n12425), .CK(clk), .Q(img[1109]), .QB(n30884) );
  DFFN img_reg_7__4__5_ ( .D(n12415), .CK(clk), .Q(img[1117]), .QB(n30821) );
  DFFN img_reg_7__2__5_ ( .D(n12399), .CK(clk), .Q(img[1133]), .QB(n30885) );
  DFFN img_reg_7__7__5_ ( .D(n12438), .CK(clk), .Q(img[1093]), .QB(n30916) );
  DFFN img_reg_7__3__5_ ( .D(n12409), .CK(clk), .Q(img[1125]), .QB(n30823) );
  DFFN img_reg_7__1__5_ ( .D(n12393), .CK(clk), .Q(img[1141]), .QB(n30940) );
  DFFN img_reg_7__0__5_ ( .D(n12383), .CK(clk), .Q(img[1149]), .QB(n30914) );
  DFFN img_reg_2__5__5_ ( .D(n11783), .CK(clk), .Q(img[1749]), .QB(n30872) );
  DFFN img_reg_2__7__5_ ( .D(n11799), .CK(clk), .Q(img[1733]), .QB(n30807) );
  DFFN img_reg_0__5__5_ ( .D(n11527), .CK(clk), .Q(img[2005]), .QB(n30891) );
  DFFN img_reg_5__5__5_ ( .D(n12169), .CK(clk), .Q(img[1365]), .QB(n30841) );
  DFFN img_reg_3__6__5_ ( .D(n11919), .CK(clk), .Q(img[1613]), .QB(n30876) );
  DFFN img_reg_3__5__5_ ( .D(n11913), .CK(clk), .Q(img[1621]), .QB(n30880) );
  DFFN img_reg_5__2__5_ ( .D(n12143), .CK(clk), .Q(img[1389]), .QB(n30842) );
  DFFN img_reg_5__4__5_ ( .D(n12159), .CK(clk), .Q(img[1373]), .QB(n30783) );
  DFFN img_reg_1__5__5_ ( .D(n11657), .CK(clk), .Q(img[1877]), .QB(n30864) );
  DFFN img_reg_5__3__5_ ( .D(n12153), .CK(clk), .Q(img[1381]), .QB(n30785) );
  DFFN img_reg_5__1__5_ ( .D(n12137), .CK(clk), .Q(img[1397]), .QB(n30952) );
  DFFN img_reg_6__4__5_ ( .D(n12289), .CK(clk), .Q(img[1245]), .QB(n30779) );
  DFFN img_reg_6__2__5_ ( .D(n12273), .CK(clk), .Q(img[1261]), .QB(n30838) );
  DFFN img_reg_6__3__5_ ( .D(n12279), .CK(clk), .Q(img[1253]), .QB(n30781) );
  DFFN img_reg_6__1__5_ ( .D(n12263), .CK(clk), .Q(img[1269]), .QB(n30949) );
  DFFN img_reg_1__6__5_ ( .D(n11663), .CK(clk), .Q(img[1869]), .QB(n30860) );
  DFFN img_reg_2__2__5_ ( .D(n11761), .CK(clk), .Q(img[1773]), .QB(n30873) );
  DFFN img_reg_14__5__4_ ( .D(n13320), .CK(clk), .Q(img[212]), .QB(n31905) );
  DFFN img_reg_12__10__4_ ( .D(n13104), .CK(clk), .Q(img[428]), .QB(n31908) );
  DFFN img_reg_15__5__4_ ( .D(n13448), .CK(clk), .Q(img[84]), .QB(n31901) );
  DFFN img_reg_14__10__4_ ( .D(n13360), .CK(clk), .Q(img[172]), .QB(n31904) );
  DFFN img_reg_1__0__5_ ( .D(n11615), .CK(clk), .Q(img[1917]), .QB(n30802) );
  DFFN img_reg_0__3__5_ ( .D(n11511), .CK(clk), .Q(img[2021]), .QB(n30831) );
  DFFN img_reg_0__2__5_ ( .D(n11505), .CK(clk), .Q(img[2029]), .QB(n30892) );
  DFFN img_reg_1__2__5_ ( .D(n11631), .CK(clk), .Q(img[1901]), .QB(n30865) );
  DFFN img_reg_2__3__5_ ( .D(n11767), .CK(clk), .Q(img[1765]), .QB(n30813) );
  DFFN img_reg_1__3__5_ ( .D(n11641), .CK(clk), .Q(img[1893]), .QB(n30805) );
  DFFN img_reg_1__1__5_ ( .D(n11625), .CK(clk), .Q(img[1909]), .QB(n30862) );
  DFFN img_reg_0__1__5_ ( .D(n11495), .CK(clk), .Q(img[2037]), .QB(n30889) );
  DFFN img_reg_3__2__5_ ( .D(n11887), .CK(clk), .Q(img[1645]), .QB(n30881) );
  DFFN img_reg_3__1__5_ ( .D(n11881), .CK(clk), .Q(img[1653]), .QB(n30878) );
  DFFN img_reg_4__5__2_ ( .D(n12042), .CK(clk), .Q(img[1490]), .QB(n30614) );
  DFFN img_reg_4__5__0_ ( .D(n12044), .CK(clk), .Q(img[1488]), .QB(n31594) );
  DFFN img_reg_4__6__2_ ( .D(n12046), .CK(clk), .Q(img[1482]), .QB(n30549) );
  DFFN img_reg_4__7__2_ ( .D(n12058), .CK(clk), .Q(img[1474]), .QB(n30661) );
  DFFN img_reg_4__6__0_ ( .D(n12052), .CK(clk), .Q(img[1480]), .QB(n31657) );
  DFFN img_reg_2__6__2_ ( .D(n11790), .CK(clk), .Q(img[1738]), .QB(n30568) );
  DFFN img_reg_0__7__2_ ( .D(n11546), .CK(clk), .Q(img[1986]), .QB(n30646) );
  DFFN img_reg_0__7__0_ ( .D(n11548), .CK(clk), .Q(img[1984]), .QB(n31558) );
  DFFN img_reg_6__5__2_ ( .D(n12298), .CK(clk), .Q(img[1234]), .QB(n30598) );
  DFFN img_reg_6__5__0_ ( .D(n12300), .CK(clk), .Q(img[1232]), .QB(n31578) );
  DFFN img_reg_3__6__2_ ( .D(n11922), .CK(clk), .Q(img[1610]), .QB(n30576) );
  DFFN img_reg_3__5__2_ ( .D(n11910), .CK(clk), .Q(img[1618]), .QB(n30572) );
  DFFN img_reg_7__6__0_ ( .D(n12436), .CK(clk), .Q(img[1096]), .QB(n31664) );
  DFFN img_reg_7__5__2_ ( .D(n12422), .CK(clk), .Q(img[1106]), .QB(n30621) );
  DFFN img_reg_7__4__2_ ( .D(n12418), .CK(clk), .Q(img[1114]), .QB(n30740) );
  DFFN img_reg_7__4__0_ ( .D(n12420), .CK(clk), .Q(img[1112]), .QB(n31697) );
  DFFN img_reg_7__2__2_ ( .D(n12402), .CK(clk), .Q(img[1130]), .QB(n30619) );
  DFFN img_reg_7__2__0_ ( .D(n12404), .CK(clk), .Q(img[1128]), .QB(n31627) );
  DFFN img_reg_7__7__2_ ( .D(n12442), .CK(clk), .Q(img[1090]), .QB(n30692) );
  DFFN img_reg_7__7__0_ ( .D(n12444), .CK(clk), .Q(img[1088]), .QB(n31550) );
  DFFN img_reg_7__3__2_ ( .D(n12406), .CK(clk), .Q(img[1122]), .QB(n30738) );
  DFFN img_reg_7__3__0_ ( .D(n12412), .CK(clk), .Q(img[1120]), .QB(n31695) );
  DFFN img_reg_7__1__0_ ( .D(n12396), .CK(clk), .Q(img[1136]), .QB(n31665) );
  DFFN img_reg_7__0__2_ ( .D(n12386), .CK(clk), .Q(img[1146]), .QB(n30694) );
  DFFN img_reg_7__0__0_ ( .D(n12388), .CK(clk), .Q(img[1144]), .QB(n31548) );
  DFFN img_reg_2__5__2_ ( .D(n11786), .CK(clk), .Q(img[1746]), .QB(n30564) );
  DFFN img_reg_2__5__0_ ( .D(n11788), .CK(clk), .Q(img[1744]), .QB(n31613) );
  DFFN img_reg_2__7__2_ ( .D(n11802), .CK(clk), .Q(img[1730]), .QB(n30680) );
  DFFN img_reg_0__6__0_ ( .D(n11540), .CK(clk), .Q(img[1992]), .QB(n31629) );
  DFFN img_reg_6__2__2_ ( .D(n12270), .CK(clk), .Q(img[1258]), .QB(n30596) );
  DFFN img_reg_1__6__2_ ( .D(n11666), .CK(clk), .Q(img[1866]), .QB(n30560) );
  DFFN img_reg_5__5__2_ ( .D(n12166), .CK(clk), .Q(img[1362]), .QB(n30602) );
  DFFN img_reg_5__5__0_ ( .D(n12172), .CK(clk), .Q(img[1360]), .QB(n31582) );
  DFFN img_reg_3__6__0_ ( .D(n11924), .CK(clk), .Q(img[1608]), .QB(n31617) );
  DFFN img_reg_3__5__0_ ( .D(n11916), .CK(clk), .Q(img[1616]), .QB(n31621) );
  DFFN img_reg_1__5__2_ ( .D(n11654), .CK(clk), .Q(img[1874]), .QB(n30556) );
  DFFN img_reg_5__2__2_ ( .D(n12146), .CK(clk), .Q(img[1386]), .QB(n30600) );
  DFFN img_reg_5__2__0_ ( .D(n12148), .CK(clk), .Q(img[1384]), .QB(n31584) );
  DFFN img_reg_5__4__2_ ( .D(n12162), .CK(clk), .Q(img[1370]), .QB(n30723) );
  DFFN img_reg_5__4__0_ ( .D(n12164), .CK(clk), .Q(img[1368]), .QB(n31678) );
  DFFN img_reg_7__6__2_ ( .D(n12434), .CK(clk), .Q(img[1098]), .QB(n30580) );
  DFFN img_reg_5__0__2_ ( .D(n12130), .CK(clk), .Q(img[1402]), .QB(n30654) );
  DFFN img_reg_1__6__0_ ( .D(n11668), .CK(clk), .Q(img[1864]), .QB(n31601) );
  DFFN img_reg_1__5__0_ ( .D(n11660), .CK(clk), .Q(img[1872]), .QB(n31605) );
  DFFN img_reg_5__3__2_ ( .D(n12150), .CK(clk), .Q(img[1378]), .QB(n30721) );
  DFFN img_reg_5__3__0_ ( .D(n12156), .CK(clk), .Q(img[1376]), .QB(n31676) );
  DFFN img_reg_5__7__2_ ( .D(n12182), .CK(clk), .Q(img[1346]), .QB(n30652) );
  DFFN img_reg_5__7__0_ ( .D(n12188), .CK(clk), .Q(img[1344]), .QB(n31520) );
  DFFN img_reg_3__7__2_ ( .D(n11926), .CK(clk), .Q(img[1602]), .QB(n30688) );
  DFFN img_reg_6__4__0_ ( .D(n12292), .CK(clk), .Q(img[1240]), .QB(n31674) );
  DFFN img_reg_0__6__2_ ( .D(n11534), .CK(clk), .Q(img[1994]), .QB(n30588) );
  DFFN img_reg_0__5__2_ ( .D(n11530), .CK(clk), .Q(img[2002]), .QB(n30584) );
  DFFN img_reg_6__4__2_ ( .D(n12286), .CK(clk), .Q(img[1242]), .QB(n30719) );
  DFFN img_reg_6__2__0_ ( .D(n12276), .CK(clk), .Q(img[1256]), .QB(n31580) );
  DFFN img_reg_6__0__2_ ( .D(n12254), .CK(clk), .Q(img[1274]), .QB(n30640) );
  DFFN img_reg_6__3__2_ ( .D(n12282), .CK(clk), .Q(img[1250]), .QB(n30717) );
  DFFN img_reg_6__7__2_ ( .D(n12314), .CK(clk), .Q(img[1218]), .QB(n30638) );
  DFFN img_reg_1__1__2_ ( .D(n11622), .CK(clk), .Q(img[1906]), .QB(n30561) );
  DFFN img_reg_2__2__2_ ( .D(n11758), .CK(clk), .Q(img[1770]), .QB(n30566) );
  DFFN img_reg_2__0__0_ ( .D(n11748), .CK(clk), .Q(img[1784]), .QB(n31536) );
  DFFN img_reg_0__1__2_ ( .D(n11498), .CK(clk), .Q(img[2034]), .QB(n30589) );
  DFFN img_reg_0__2__0_ ( .D(n11508), .CK(clk), .Q(img[2024]), .QB(n31635) );
  DFFN img_reg_2__2__0_ ( .D(n11764), .CK(clk), .Q(img[1768]), .QB(n31615) );
  DFFN img_reg_1__2__0_ ( .D(n11636), .CK(clk), .Q(img[1896]), .QB(n31607) );
  DFFN img_reg_3__3__0_ ( .D(n11900), .CK(clk), .Q(img[1632]), .QB(n31542) );
  DFFN img_reg_2__3__0_ ( .D(n11772), .CK(clk), .Q(img[1760]), .QB(n31534) );
  DFFN img_reg_2__1__2_ ( .D(n11754), .CK(clk), .Q(img[1778]), .QB(n30569) );
  DFFN img_reg_2__1__0_ ( .D(n11756), .CK(clk), .Q(img[1776]), .QB(n31611) );
  DFFN img_reg_3__2__0_ ( .D(n11892), .CK(clk), .Q(img[1640]), .QB(n31623) );
  DFFN img_reg_3__1__0_ ( .D(n11884), .CK(clk), .Q(img[1648]), .QB(n31619) );
  DFFN img_reg_3__0__0_ ( .D(n11876), .CK(clk), .Q(img[1656]), .QB(n31544) );
  DFFN img_reg_2__0__2_ ( .D(n11742), .CK(clk), .Q(img[1786]), .QB(n30682) );
  DFFN img_reg_3__3__2_ ( .D(n11893), .CK(clk), .Q(img[1634]), .QB(n30686) );
  DFFN img_reg_1__1__0_ ( .D(n11628), .CK(clk), .Q(img[1904]), .QB(n31603) );
  DFFN img_reg_0__3__2_ ( .D(n11514), .CK(clk), .Q(img[2018]), .QB(n30644) );
  DFFN img_reg_0__3__0_ ( .D(n11516), .CK(clk), .Q(img[2016]), .QB(n31554) );
  DFFN img_reg_0__1__0_ ( .D(n11500), .CK(clk), .Q(img[2032]), .QB(n31631) );
  DFFN img_reg_3__2__2_ ( .D(n11890), .CK(clk), .Q(img[1642]), .QB(n30574) );
  DFFN img_reg_3__1__2_ ( .D(n11878), .CK(clk), .Q(img[1650]), .QB(n30577) );
  DFFN img_reg_6__6__3_ ( .D(n12303), .CK(clk), .Q(img[1227]), .QB(n31394) );
  DFFN img_reg_6__5__3_ ( .D(n12297), .CK(clk), .Q(img[1235]), .QB(n31263) );
  DFFN img_reg_4__7__3_ ( .D(n12057), .CK(clk), .Q(img[1475]), .QB(n31355) );
  DFFN img_reg_0__7__3_ ( .D(n11545), .CK(clk), .Q(img[1987]), .QB(n31388) );
  DFFN img_reg_5__6__3_ ( .D(n12177), .CK(clk), .Q(img[1355]), .QB(n31398) );
  DFFN img_reg_3__6__3_ ( .D(n11921), .CK(clk), .Q(img[1611]), .QB(n31298) );
  DFFN img_reg_1__5__3_ ( .D(n11655), .CK(clk), .Q(img[1875]), .QB(n31288) );
  DFFN img_reg_2__5__3_ ( .D(n11785), .CK(clk), .Q(img[1747]), .QB(n31294) );
  DFFN img_reg_0__6__3_ ( .D(n11535), .CK(clk), .Q(img[1995]), .QB(n31310) );
  DFFN img_reg_0__5__3_ ( .D(n11529), .CK(clk), .Q(img[2003]), .QB(n31314) );
  DFFN img_reg_6__2__3_ ( .D(n12271), .CK(clk), .Q(img[1259]), .QB(n31264) );
  DFFN img_reg_6__0__3_ ( .D(n12255), .CK(clk), .Q(img[1275]), .QB(n31337) );
  DFFN img_reg_5__2__3_ ( .D(n12145), .CK(clk), .Q(img[1387]), .QB(n31268) );
  DFFN img_reg_5__0__3_ ( .D(n12129), .CK(clk), .Q(img[1403]), .QB(n31341) );
  DFFN img_reg_6__4__3_ ( .D(n12287), .CK(clk), .Q(img[1243]), .QB(n31447) );
  DFFN img_reg_6__3__3_ ( .D(n12281), .CK(clk), .Q(img[1251]), .QB(n31445) );
  DFFN img_reg_6__1__3_ ( .D(n12265), .CK(clk), .Q(img[1267]), .QB(n31395) );
  DFFN img_reg_5__4__3_ ( .D(n12161), .CK(clk), .Q(img[1371]), .QB(n31451) );
  DFFN img_reg_5__3__3_ ( .D(n12151), .CK(clk), .Q(img[1379]), .QB(n31449) );
  DFFN img_reg_7__6__3_ ( .D(n12433), .CK(clk), .Q(img[1099]), .QB(n31416) );
  DFFN img_reg_7__5__3_ ( .D(n12423), .CK(clk), .Q(img[1107]), .QB(n31306) );
  DFFN img_reg_7__4__3_ ( .D(n12417), .CK(clk), .Q(img[1115]), .QB(n31440) );
  DFFN img_reg_7__3__3_ ( .D(n12407), .CK(clk), .Q(img[1123]), .QB(n31438) );
  DFFN img_reg_7__2__3_ ( .D(n12401), .CK(clk), .Q(img[1131]), .QB(n31307) );
  DFFN img_reg_7__1__3_ ( .D(n12391), .CK(clk), .Q(img[1139]), .QB(n31417) );
  DFFN img_reg_6__7__3_ ( .D(n12313), .CK(clk), .Q(img[1219]), .QB(n31339) );
  DFFN img_reg_5__7__3_ ( .D(n12183), .CK(clk), .Q(img[1347]), .QB(n31343) );
  DFFN img_reg_3__7__3_ ( .D(n11927), .CK(clk), .Q(img[1603]), .QB(n31380) );
  DFFN img_reg_2__7__3_ ( .D(n11801), .CK(clk), .Q(img[1731]), .QB(n31373) );
  DFFN img_reg_1__7__3_ ( .D(n11671), .CK(clk), .Q(img[1859]), .QB(n31365) );
  DFFN img_reg_0__1__3_ ( .D(n11497), .CK(clk), .Q(img[2035]), .QB(n31312) );
  DFFN img_reg_2__0__3_ ( .D(n11743), .CK(clk), .Q(img[1787]), .QB(n31371) );
  DFFN img_reg_1__3__3_ ( .D(n11639), .CK(clk), .Q(img[1891]), .QB(n31361) );
  DFFN img_reg_3__3__3_ ( .D(n11894), .CK(clk), .Q(img[1635]), .QB(n31376) );
  DFFN img_reg_2__3__3_ ( .D(n11769), .CK(clk), .Q(img[1763]), .QB(n31369) );
  DFFN img_reg_2__1__3_ ( .D(n11753), .CK(clk), .Q(img[1779]), .QB(n31292) );
  DFFN img_reg_3__2__3_ ( .D(n11889), .CK(clk), .Q(img[1643]), .QB(n31303) );
  DFFN img_reg_3__1__3_ ( .D(n11879), .CK(clk), .Q(img[1651]), .QB(n31300) );
  DFFN img_reg_3__0__3_ ( .D(n11873), .CK(clk), .Q(img[1659]), .QB(n31378) );
  DFFN img_reg_4__6__6_ ( .D(n12050), .CK(clk), .Q(img[1486]), .QB(n30365) );
  DFFN img_reg_4__6__1_ ( .D(n12045), .CK(clk), .Q(img[1481]), .QB(n31202) );
  DFFN img_reg_2__6__6_ ( .D(n11794), .CK(clk), .Q(img[1742]), .QB(n30384) );
  DFFN img_reg_4__7__1_ ( .D(n12059), .CK(clk), .Q(img[1473]), .QB(n31031) );
  DFFN img_reg_6__6__1_ ( .D(n12301), .CK(clk), .Q(img[1225]), .QB(n31183) );
  DFFN img_reg_2__6__1_ ( .D(n11789), .CK(clk), .Q(img[1737]), .QB(n31155) );
  DFFN img_reg_0__7__6_ ( .D(n11542), .CK(clk), .Q(img[1990]), .QB(n30343) );
  DFFN img_reg_0__7__1_ ( .D(n11547), .CK(clk), .Q(img[1985]), .QB(n31071) );
  DFFN img_reg_6__6__6_ ( .D(n12306), .CK(clk), .Q(img[1230]), .QB(n30349) );
  DFFN img_reg_3__6__1_ ( .D(n11923), .CK(clk), .Q(img[1609]), .QB(n31163) );
  DFFN img_reg_3__5__6_ ( .D(n11914), .CK(clk), .Q(img[1622]), .QB(n30388) );
  DFFN img_reg_3__5__1_ ( .D(n11909), .CK(clk), .Q(img[1617]), .QB(n31169) );
  DFFN img_reg_1__6__1_ ( .D(n11667), .CK(clk), .Q(img[1865]), .QB(n31147) );
  DFFN img_reg_7__6__6_ ( .D(n12430), .CK(clk), .Q(img[1102]), .QB(n30396) );
  DFFN img_reg_7__6__1_ ( .D(n12435), .CK(clk), .Q(img[1097]), .QB(n31208) );
  DFFN img_reg_7__4__6_ ( .D(n12414), .CK(clk), .Q(img[1118]), .QB(n30435) );
  DFFN img_reg_7__4__1_ ( .D(n12419), .CK(clk), .Q(img[1113]), .QB(n31102) );
  DFFN img_reg_7__2__6_ ( .D(n12398), .CK(clk), .Q(img[1134]), .QB(n30491) );
  DFFN img_reg_7__2__1_ ( .D(n12403), .CK(clk), .Q(img[1129]), .QB(n31171) );
  DFFN img_reg_7__7__6_ ( .D(n12439), .CK(clk), .Q(img[1094]), .QB(n30335) );
  DFFN img_reg_7__7__1_ ( .D(n12443), .CK(clk), .Q(img[1089]), .QB(n31063) );
  DFFN img_reg_7__3__6_ ( .D(n12410), .CK(clk), .Q(img[1126]), .QB(n30436) );
  DFFN img_reg_7__1__6_ ( .D(n12394), .CK(clk), .Q(img[1142]), .QB(n30398) );
  DFFN img_reg_7__1__1_ ( .D(n12389), .CK(clk), .Q(img[1137]), .QB(n31210) );
  DFFN img_reg_7__0__6_ ( .D(n12382), .CK(clk), .Q(img[1150]), .QB(n30333) );
  DFFN img_reg_2__5__6_ ( .D(n11782), .CK(clk), .Q(img[1750]), .QB(n30380) );
  DFFN img_reg_0__5__1_ ( .D(n11531), .CK(clk), .Q(img[2001]), .QB(n31181) );
  DFFN img_reg_2__7__6_ ( .D(n11798), .CK(clk), .Q(img[1734]), .QB(n30323) );
  DFFN img_reg_1__6__6_ ( .D(n11662), .CK(clk), .Q(img[1870]), .QB(n30376) );
  DFFN img_reg_1__5__6_ ( .D(n11658), .CK(clk), .Q(img[1878]), .QB(n30372) );
  DFFN img_reg_1__5__1_ ( .D(n11653), .CK(clk), .Q(img[1873]), .QB(n31153) );
  DFFN img_reg_6__1__6_ ( .D(n12262), .CK(clk), .Q(img[1270]), .QB(n30351) );
  DFFN img_reg_5__6__6_ ( .D(n12174), .CK(clk), .Q(img[1358]), .QB(n30353) );
  DFFN img_reg_5__6__1_ ( .D(n12179), .CK(clk), .Q(img[1353]), .QB(n31192) );
  DFFN img_reg_5__5__6_ ( .D(n12170), .CK(clk), .Q(img[1366]), .QB(n30484) );
  DFFN img_reg_5__5__1_ ( .D(n12165), .CK(clk), .Q(img[1361]), .QB(n31130) );
  DFFN img_reg_5__4__1_ ( .D(n12163), .CK(clk), .Q(img[1369]), .QB(n31083) );
  DFFN img_reg_7__5__6_ ( .D(n12426), .CK(clk), .Q(img[1110]), .QB(n30492) );
  DFFN img_reg_7__5__1_ ( .D(n12421), .CK(clk), .Q(img[1105]), .QB(n31173) );
  DFFN img_reg_5__0__6_ ( .D(n12126), .CK(clk), .Q(img[1406]), .QB(n30291) );
  DFFN img_reg_5__0__1_ ( .D(n12131), .CK(clk), .Q(img[1401]), .QB(n31021) );
  DFFN img_reg_5__3__1_ ( .D(n12149), .CK(clk), .Q(img[1377]), .QB(n31082) );
  DFFN img_reg_5__1__6_ ( .D(n12138), .CK(clk), .Q(img[1398]), .QB(n30355) );
  DFFN img_reg_5__7__6_ ( .D(n12186), .CK(clk), .Q(img[1350]), .QB(n30293) );
  DFFN img_reg_5__7__1_ ( .D(n12181), .CK(clk), .Q(img[1345]), .QB(n31020) );
  DFFN img_reg_3__7__6_ ( .D(n11930), .CK(clk), .Q(img[1606]), .QB(n30331) );
  DFFN img_reg_3__7__1_ ( .D(n11925), .CK(clk), .Q(img[1601]), .QB(n31059) );
  DFFN img_reg_2__5__1_ ( .D(n11787), .CK(clk), .Q(img[1745]), .QB(n31161) );
  DFFN img_reg_1__7__6_ ( .D(n11674), .CK(clk), .Q(img[1862]), .QB(n30315) );
  DFFN img_reg_1__7__1_ ( .D(n11669), .CK(clk), .Q(img[1857]), .QB(n31043) );
  DFFN img_reg_0__5__6_ ( .D(n11526), .CK(clk), .Q(img[2006]), .QB(n30400) );
  DFFN img_reg_6__4__6_ ( .D(n12290), .CK(clk), .Q(img[1246]), .QB(n30412) );
  DFFN img_reg_6__4__1_ ( .D(n12285), .CK(clk), .Q(img[1241]), .QB(n31079) );
  DFFN img_reg_6__0__6_ ( .D(n12258), .CK(clk), .Q(img[1278]), .QB(n30287) );
  DFFN img_reg_6__0__1_ ( .D(n12253), .CK(clk), .Q(img[1273]), .QB(n31017) );
  DFFN img_reg_6__3__1_ ( .D(n12283), .CK(clk), .Q(img[1249]), .QB(n31078) );
  DFFN img_reg_6__1__1_ ( .D(n12267), .CK(clk), .Q(img[1265]), .QB(n31185) );
  DFFN img_reg_6__7__6_ ( .D(n12310), .CK(clk), .Q(img[1222]), .QB(n30289) );
  DFFN img_reg_6__7__1_ ( .D(n12315), .CK(clk), .Q(img[1217]), .QB(n31016) );
  DFFN img_reg_5__1__1_ ( .D(n12133), .CK(clk), .Q(img[1393]), .QB(n31194) );
  DFFN img_reg_3__0__6_ ( .D(n11870), .CK(clk), .Q(img[1662]), .QB(n30329) );
  DFFN img_reg_4__6__7_ ( .D(n12051), .CK(clk), .Q(img[1487]), .QB(n30061) );
  DFFN img_reg_6__5__7_ ( .D(n12293), .CK(clk), .Q(img[1239]), .QB(n30199) );
  DFFN img_reg_4__7__7_ ( .D(n12053), .CK(clk), .Q(img[1479]), .QB(n30187) );
  DFFN img_reg_6__6__7_ ( .D(n12307), .CK(clk), .Q(img[1231]), .QB(n30045) );
  DFFN img_reg_7__6__7_ ( .D(n12429), .CK(clk), .Q(img[1103]), .QB(n30092) );
  DFFN img_reg_7__5__7_ ( .D(n12427), .CK(clk), .Q(img[1111]), .QB(n30222) );
  DFFN img_reg_7__2__7_ ( .D(n12397), .CK(clk), .Q(img[1135]), .QB(n30223) );
  DFFN img_reg_7__7__7_ ( .D(n12440), .CK(clk), .Q(img[1095]), .QB(n30193) );
  DFFN img_reg_7__3__7_ ( .D(n12411), .CK(clk), .Q(img[1127]), .QB(n30154) );
  DFFN img_reg_7__1__7_ ( .D(n12395), .CK(clk), .Q(img[1143]), .QB(n30090) );
  DFFN img_reg_7__0__7_ ( .D(n12381), .CK(clk), .Q(img[1151]), .QB(n30191) );
  DFFN img_reg_2__7__7_ ( .D(n11797), .CK(clk), .Q(img[1735]), .QB(n30137) );
  DFFN img_reg_1__5__7_ ( .D(n11659), .CK(clk), .Q(img[1879]), .QB(n30066) );
  DFFN img_reg_0__6__7_ ( .D(n11539), .CK(clk), .Q(img[1999]), .QB(n30100) );
  DFFN img_reg_5__6__7_ ( .D(n12173), .CK(clk), .Q(img[1359]), .QB(n30049) );
  DFFN img_reg_5__5__7_ ( .D(n12171), .CK(clk), .Q(img[1367]), .QB(n30203) );
  DFFN img_reg_3__6__7_ ( .D(n11917), .CK(clk), .Q(img[1615]), .QB(n30088) );
  DFFN img_reg_5__0__7_ ( .D(n12125), .CK(clk), .Q(img[1407]), .QB(n30173) );
  DFFN img_reg_5__3__7_ ( .D(n12155), .CK(clk), .Q(img[1383]), .QB(n30111) );
  DFFN img_reg_5__1__7_ ( .D(n12139), .CK(clk), .Q(img[1399]), .QB(n30047) );
  DFFN img_reg_5__7__7_ ( .D(n12187), .CK(clk), .Q(img[1351]), .QB(n30175) );
  DFFN img_reg_3__7__7_ ( .D(n11931), .CK(clk), .Q(img[1607]), .QB(n30145) );
  DFFN img_reg_2__5__7_ ( .D(n11781), .CK(clk), .Q(img[1751]), .QB(n30074) );
  DFFN img_reg_1__7__7_ ( .D(n11675), .CK(clk), .Q(img[1863]), .QB(n30129) );
  DFFN img_reg_0__5__7_ ( .D(n11525), .CK(clk), .Q(img[2007]), .QB(n30094) );
  DFFN img_reg_6__4__7_ ( .D(n12291), .CK(clk), .Q(img[1247]), .QB(n30106) );
  DFFN img_reg_6__2__7_ ( .D(n12275), .CK(clk), .Q(img[1263]), .QB(n30200) );
  DFFN img_reg_6__0__7_ ( .D(n12259), .CK(clk), .Q(img[1279]), .QB(n30169) );
  DFFN img_reg_6__3__7_ ( .D(n12277), .CK(clk), .Q(img[1255]), .QB(n30107) );
  DFFN img_reg_6__1__7_ ( .D(n12261), .CK(clk), .Q(img[1271]), .QB(n30043) );
  DFFN img_reg_6__7__7_ ( .D(n12309), .CK(clk), .Q(img[1223]), .QB(n30171) );
  DFFN img_reg_2__2__6_ ( .D(n11762), .CK(clk), .Q(img[1774]), .QB(n30382) );
  DFFN img_reg_0__2__6_ ( .D(n11506), .CK(clk), .Q(img[2030]), .QB(n30402) );
  DFFN img_reg_0__2__1_ ( .D(n11501), .CK(clk), .Q(img[2025]), .QB(n31179) );
  DFFN img_reg_1__2__1_ ( .D(n11635), .CK(clk), .Q(img[1897]), .QB(n31151) );
  DFFN img_reg_3__3__1_ ( .D(n11899), .CK(clk), .Q(img[1633]), .QB(n31057) );
  DFFN img_reg_2__1__1_ ( .D(n11755), .CK(clk), .Q(img[1777]), .QB(n31157) );
  DFFN img_reg_1__1__1_ ( .D(n11621), .CK(clk), .Q(img[1905]), .QB(n31149) );
  DFFN img_reg_0__3__1_ ( .D(n11515), .CK(clk), .Q(img[2017]), .QB(n31069) );
  DFFN img_reg_3__1__1_ ( .D(n11877), .CK(clk), .Q(img[1649]), .QB(n31165) );
  DFFN img_reg_2__0__6_ ( .D(n11746), .CK(clk), .Q(img[1790]), .QB(n30321) );
  DFFN img_reg_1__2__6_ ( .D(n11630), .CK(clk), .Q(img[1902]), .QB(n30374) );
  DFFN img_reg_3__3__6_ ( .D(n11897), .CK(clk), .Q(img[1638]), .QB(n30327) );
  DFFN img_reg_2__3__6_ ( .D(n11766), .CK(clk), .Q(img[1766]), .QB(n30319) );
  DFFN img_reg_2__1__6_ ( .D(n11750), .CK(clk), .Q(img[1782]), .QB(n30386) );
  DFFN img_reg_0__1__1_ ( .D(n11499), .CK(clk), .Q(img[2033]), .QB(n31177) );
  DFFN img_reg_3__2__6_ ( .D(n11886), .CK(clk), .Q(img[1646]), .QB(n30390) );
  DFFN img_reg_3__2__1_ ( .D(n11891), .CK(clk), .Q(img[1641]), .QB(n31167) );
  DFFN img_reg_3__1__6_ ( .D(n11882), .CK(clk), .Q(img[1654]), .QB(n30394) );
  DFFN img_reg_0__2__7_ ( .D(n11507), .CK(clk), .Q(img[2031]), .QB(n30096) );
  DFFN img_reg_0__3__7_ ( .D(n11509), .CK(clk), .Q(img[2023]), .QB(n30162) );
  DFFN img_reg_2__0__7_ ( .D(n11747), .CK(clk), .Q(img[1791]), .QB(n30139) );
  DFFN img_reg_1__2__7_ ( .D(n11629), .CK(clk), .Q(img[1903]), .QB(n30068) );
  DFFN img_reg_1__0__7_ ( .D(n11613), .CK(clk), .Q(img[1919]), .QB(n30131) );
  DFFN img_reg_2__3__7_ ( .D(n11765), .CK(clk), .Q(img[1767]), .QB(n30142) );
  DFFN img_reg_1__3__7_ ( .D(n11643), .CK(clk), .Q(img[1895]), .QB(n30134) );
  DFFN img_reg_3__2__7_ ( .D(n11885), .CK(clk), .Q(img[1647]), .QB(n30084) );
  DFFN img_reg_3__0__7_ ( .D(n11869), .CK(clk), .Q(img[1663]), .QB(n30147) );
  DFFN img_reg_4__5__4_ ( .D(n12040), .CK(clk), .Q(img[1492]), .QB(n31888) );
  DFFN img_reg_4__7__4_ ( .D(n12056), .CK(clk), .Q(img[1476]), .QB(n31827) );
  DFFN img_reg_6__6__4_ ( .D(n12304), .CK(clk), .Q(img[1228]), .QB(n31749) );
  DFFN img_reg_6__5__4_ ( .D(n12296), .CK(clk), .Q(img[1236]), .QB(n31872) );
  DFFN img_reg_7__6__4_ ( .D(n12432), .CK(clk), .Q(img[1100]), .QB(n31796) );
  DFFN img_reg_7__5__4_ ( .D(n12424), .CK(clk), .Q(img[1108]), .QB(n31895) );
  DFFN img_reg_7__4__4_ ( .D(n12416), .CK(clk), .Q(img[1116]), .QB(n31916) );
  DFFN img_reg_7__2__4_ ( .D(n12400), .CK(clk), .Q(img[1132]), .QB(n31897) );
  DFFN img_reg_5__3__4_ ( .D(n12152), .CK(clk), .Q(img[1380]), .QB(n31932) );
  DFFN img_reg_7__7__4_ ( .D(n12437), .CK(clk), .Q(img[1092]), .QB(n31857) );
  DFFN img_reg_7__0__4_ ( .D(n12384), .CK(clk), .Q(img[1148]), .QB(n31856) );
  DFFN img_reg_2__5__4_ ( .D(n11784), .CK(clk), .Q(img[1748]), .QB(n31778) );
  DFFN img_reg_6__2__4_ ( .D(n12272), .CK(clk), .Q(img[1260]), .QB(n31874) );
  DFFN img_reg_1__6__4_ ( .D(n11664), .CK(clk), .Q(img[1868]), .QB(n31776) );
  DFFN img_reg_0__6__4_ ( .D(n11536), .CK(clk), .Q(img[1996]), .QB(n31804) );
  DFFN img_reg_5__6__4_ ( .D(n12176), .CK(clk), .Q(img[1356]), .QB(n31753) );
  DFFN img_reg_5__5__4_ ( .D(n12168), .CK(clk), .Q(img[1364]), .QB(n31876) );
  DFFN img_reg_3__5__4_ ( .D(n11912), .CK(clk), .Q(img[1620]), .QB(n31786) );
  DFFN img_reg_5__2__4_ ( .D(n12144), .CK(clk), .Q(img[1388]), .QB(n31878) );
  DFFN img_reg_5__4__4_ ( .D(n12160), .CK(clk), .Q(img[1372]), .QB(n31930) );
  DFFN img_reg_1__5__4_ ( .D(n11656), .CK(clk), .Q(img[1876]), .QB(n31770) );
  DFFN img_reg_5__1__4_ ( .D(n12136), .CK(clk), .Q(img[1396]), .QB(n31751) );
  DFFN img_reg_1__7__4_ ( .D(n11672), .CK(clk), .Q(img[1860]), .QB(n31837) );
  DFFN img_reg_6__4__4_ ( .D(n12288), .CK(clk), .Q(img[1244]), .QB(n31922) );
  DFFN img_reg_6__0__4_ ( .D(n12256), .CK(clk), .Q(img[1276]), .QB(n31810) );
  DFFN img_reg_6__1__4_ ( .D(n12264), .CK(clk), .Q(img[1268]), .QB(n31747) );
  DFFN img_reg_6__7__4_ ( .D(n12312), .CK(clk), .Q(img[1220]), .QB(n31811) );
  DFFN img_reg_5__7__4_ ( .D(n12184), .CK(clk), .Q(img[1348]), .QB(n31815) );
  DFFN img_reg_1__0__4_ ( .D(n11616), .CK(clk), .Q(img[1916]), .QB(n31836) );
  DFFN img_reg_2__1__4_ ( .D(n11752), .CK(clk), .Q(img[1780]), .QB(n31782) );
  DFFN img_reg_1__1__4_ ( .D(n11624), .CK(clk), .Q(img[1908]), .QB(n31774) );
  DFFN img_reg_0__3__4_ ( .D(n11512), .CK(clk), .Q(img[2020]), .QB(n31862) );
  DFFN img_reg_3__1__4_ ( .D(n11880), .CK(clk), .Q(img[1652]), .QB(n31790) );
  DFFN img_reg_2__0__4_ ( .D(n11744), .CK(clk), .Q(img[1788]), .QB(n31844) );
  DFFN img_reg_1__2__4_ ( .D(n11632), .CK(clk), .Q(img[1900]), .QB(n31772) );
  DFFN img_reg_1__3__4_ ( .D(n11640), .CK(clk), .Q(img[1892]), .QB(n31834) );
  DFFN img_reg_0__1__4_ ( .D(n11496), .CK(clk), .Q(img[2036]), .QB(n31802) );
  DFFN img_reg_3__0__4_ ( .D(n11872), .CK(clk), .Q(img[1660]), .QB(n31852) );
  DFFN img_reg_0__13__5_ ( .D(n11591), .CK(clk), .Q(img[1941]), .QB(n30893) );
  DFFN img_reg_14__8__5_ ( .D(n13345), .CK(clk), .Q(img[189]), .QB(n30894) );
  DFFN img_reg_14__7__5_ ( .D(n13335), .CK(clk), .Q(img[197]), .QB(n30895) );
  DFFN img_reg_12__8__5_ ( .D(n13090), .CK(clk), .Q(img[445]), .QB(n30906) );
  DFFN img_reg_12__7__5_ ( .D(n13079), .CK(clk), .Q(img[453]), .QB(n30907) );
  DFFN img_reg_15__7__5_ ( .D(n13465), .CK(clk), .Q(img[69]), .QB(n30897) );
  DFFN img_reg_6__8__5_ ( .D(n12321), .CK(clk), .Q(img[1213]), .QB(n30899) );
  DFFN img_reg_5__9__3_ ( .D(n12199), .CK(clk), .Q(img[1331]), .QB(n31397) );
  DFFN img_reg_8__7__5_ ( .D(n12567), .CK(clk), .Q(img[965]), .QB(n30903) );
  DFFN img_reg_2__12__3_ ( .D(n11839), .CK(clk), .Q(img[1691]), .QB(n31368) );
  DFFN img_reg_0__12__3_ ( .D(n11583), .CK(clk), .Q(img[1947]), .QB(n31384) );
  DFFN img_reg_0__8__3_ ( .D(n11551), .CK(clk), .Q(img[1979]), .QB(n31387) );
  DFFN img_reg_3__12__3_ ( .D(n11969), .CK(clk), .Q(img[1563]), .QB(n31375) );
  DFFN img_reg_15__1__3_ ( .D(n13415), .CK(clk), .Q(img[115]), .QB(n31391) );
  DFFN img_reg_7__10__0_ ( .D(n12468), .CK(clk), .Q(img[1064]), .QB(n31624) );
  DFFN img_reg_2__9__0_ ( .D(n11820), .CK(clk), .Q(img[1712]), .QB(n31608) );
  DFFN img_reg_3__10__0_ ( .D(n11956), .CK(clk), .Q(img[1576]), .QB(n31620) );
  DFFN img_reg_14__15__2_ ( .D(n13402), .CK(clk), .Q(img[130]), .QB(n30655) );
  DFFN img_reg_7__13__0_ ( .D(n12492), .CK(clk), .Q(img[1040]), .QB(n31626) );
  DFFN img_reg_2__13__0_ ( .D(n11852), .CK(clk), .Q(img[1680]), .QB(n31614) );
  DFFN img_reg_0__13__0_ ( .D(n11596), .CK(clk), .Q(img[1936]), .QB(n31634) );
  DFFN img_reg_5__9__0_ ( .D(n12204), .CK(clk), .Q(img[1328]), .QB(n31644) );
  DFFN img_reg_2__14__0_ ( .D(n11860), .CK(clk), .Q(img[1672]), .QB(n31610) );
  DFFN img_reg_0__14__0_ ( .D(n11604), .CK(clk), .Q(img[1928]), .QB(n31630) );
  DFFN img_reg_14__0__2_ ( .D(n13277), .CK(clk), .Q(img[250]), .QB(n30656) );
  DFFN img_reg_1__8__2_ ( .D(n11682), .CK(clk), .Q(img[1850]), .QB(n30671) );
  DFFN img_reg_15__1__0_ ( .D(n13420), .CK(clk), .Q(img[112]), .QB(n31638) );
  DFFN img_reg_7__10__5_ ( .D(n12463), .CK(clk), .Q(img[1069]), .QB(n30883) );
  DFFN img_reg_2__9__5_ ( .D(n11815), .CK(clk), .Q(img[1717]), .QB(n30867) );
  DFFN img_reg_5__11__5_ ( .D(n12217), .CK(clk), .Q(img[1317]), .QB(n30782) );
  DFFN img_reg_3__10__5_ ( .D(n11951), .CK(clk), .Q(img[1581]), .QB(n30879) );
  DFFN img_reg_1__10__5_ ( .D(n11695), .CK(clk), .Q(img[1837]), .QB(n30863) );
  DFFN img_reg_4__12__5_ ( .D(n12097), .CK(clk), .Q(img[1437]), .QB(n30796) );
  DFFN img_reg_6__11__5_ ( .D(n12343), .CK(clk), .Q(img[1189]), .QB(n30778) );
  DFFN img_reg_7__13__5_ ( .D(n12488), .CK(clk), .Q(img[1045]), .QB(n30886) );
  DFFN img_reg_5__13__5_ ( .D(n12233), .CK(clk), .Q(img[1301]), .QB(n30843) );
  DFFN img_reg_3__13__5_ ( .D(n11977), .CK(clk), .Q(img[1557]), .QB(n30882) );
  DFFN img_reg_2__13__5_ ( .D(n11847), .CK(clk), .Q(img[1685]), .QB(n30874) );
  DFFN img_reg_1__13__5_ ( .D(n11721), .CK(clk), .Q(img[1813]), .QB(n30866) );
  DFFN img_reg_7__9__5_ ( .D(n12457), .CK(clk), .Q(img[1077]), .QB(n30941) );
  DFFN img_reg_5__9__5_ ( .D(n12201), .CK(clk), .Q(img[1333]), .QB(n30953) );
  DFFN img_reg_1__9__5_ ( .D(n11689), .CK(clk), .Q(img[1845]), .QB(n30859) );
  DFFN img_reg_14__11__5_ ( .D(n13367), .CK(clk), .Q(img[165]), .QB(n31001) );
  DFFN img_reg_14__9__5_ ( .D(n13351), .CK(clk), .Q(img[181]), .QB(n30957) );
  DFFN img_reg_14__2__5_ ( .D(n13297), .CK(clk), .Q(img[237]), .QB(n30846) );
  DFFN img_reg_2__14__5_ ( .D(n11857), .CK(clk), .Q(img[1677]), .QB(n30869) );
  DFFN img_reg_0__14__5_ ( .D(n11601), .CK(clk), .Q(img[1933]), .QB(n30888) );
  DFFN img_reg_2__12__5_ ( .D(n11841), .CK(clk), .Q(img[1693]), .QB(n30812) );
  DFFN img_reg_0__12__5_ ( .D(n11585), .CK(clk), .Q(img[1949]), .QB(n30830) );
  DFFN img_reg_14__13__5_ ( .D(n13383), .CK(clk), .Q(img[149]), .QB(n30847) );
  DFFN img_reg_14__6__5_ ( .D(n13329), .CK(clk), .Q(img[205]), .QB(n30958) );
  DFFN img_reg_14__12__5_ ( .D(n13377), .CK(clk), .Q(img[157]), .QB(n30788) );
  DFFN img_reg_12__11__5_ ( .D(n13111), .CK(clk), .Q(img[421]), .QB(n31005) );
  DFFN img_reg_14__3__5_ ( .D(n13303), .CK(clk), .Q(img[229]), .QB(n30789) );
  DFFN img_reg_14__1__5_ ( .D(n13287), .CK(clk), .Q(img[245]), .QB(n30976) );
  DFFN img_reg_14__0__5_ ( .D(n13280), .CK(clk), .Q(img[253]), .QB(n30983) );
  DFFN img_reg_12__3__5_ ( .D(n13047), .CK(clk), .Q(img[485]), .QB(n30793) );
  DFFN img_reg_12__2__5_ ( .D(n13041), .CK(clk), .Q(img[493]), .QB(n30850) );
  DFFN img_reg_12__1__5_ ( .D(n13031), .CK(clk), .Q(img[501]), .QB(n30968) );
  DFFN img_reg_14__4__5_ ( .D(n13313), .CK(clk), .Q(img[221]), .QB(n31002) );
  DFFN img_reg_12__4__5_ ( .D(n13057), .CK(clk), .Q(img[477]), .QB(n31006) );
  DFFN img_reg_0__8__5_ ( .D(n11553), .CK(clk), .Q(img[1981]), .QB(n30824) );
  DFFN img_reg_15__12__5_ ( .D(n13503), .CK(clk), .Q(img[29]), .QB(n30776) );
  DFFN img_reg_15__11__5_ ( .D(n13497), .CK(clk), .Q(img[37]), .QB(n30997) );
  DFFN img_reg_15__5__5_ ( .D(n13449), .CK(clk), .Q(img[85]), .QB(n30924) );
  DFFN img_reg_12__12__5_ ( .D(n13121), .CK(clk), .Q(img[413]), .QB(n30792) );
  DFFN img_reg_3__12__5_ ( .D(n11967), .CK(clk), .Q(img[1565]), .QB(n30819) );
  DFFN img_reg_1__12__5_ ( .D(n11711), .CK(clk), .Q(img[1821]), .QB(n30804) );
  DFFN img_reg_15__4__5_ ( .D(n13439), .CK(clk), .Q(img[93]), .QB(n30998) );
  DFFN img_reg_15__3__5_ ( .D(n13433), .CK(clk), .Q(img[101]), .QB(n30777) );
  DFFN img_reg_15__1__5_ ( .D(n13417), .CK(clk), .Q(img[117]), .QB(n30970) );
  DFFN img_reg_15__0__5_ ( .D(n13407), .CK(clk), .Q(img[125]), .QB(n30989) );
  DFFN img_reg_15__2__5_ ( .D(n13423), .CK(clk), .Q(img[109]), .QB(n30834) );
  DFFN img_reg_11__12__5_ ( .D(n12991), .CK(clk), .Q(img[541]), .QB(n30774) );
  DFFN img_reg_10__12__5_ ( .D(n12865), .CK(clk), .Q(img[669]), .QB(n30798) );
  DFFN img_reg_8__12__5_ ( .D(n12609), .CK(clk), .Q(img[925]), .QB(n30786) );
  DFFN img_reg_6__12__5_ ( .D(n12353), .CK(clk), .Q(img[1181]), .QB(n30780) );
  DFFN img_reg_8__5__5_ ( .D(n12551), .CK(clk), .Q(img[981]), .QB(n30926) );
  DFFN img_reg_8__4__5_ ( .D(n12545), .CK(clk), .Q(img[989]), .QB(n31000) );
  DFFN img_reg_8__3__5_ ( .D(n12535), .CK(clk), .Q(img[997]), .QB(n30787) );
  DFFN img_reg_8__2__5_ ( .D(n12529), .CK(clk), .Q(img[1005]), .QB(n30844) );
  DFFN img_reg_8__1__5_ ( .D(n12519), .CK(clk), .Q(img[1013]), .QB(n30974) );
  DFFN img_reg_11__10__5_ ( .D(n12975), .CK(clk), .Q(img[557]), .QB(n30921) );
  DFFN img_reg_11__8__5_ ( .D(n12959), .CK(clk), .Q(img[573]), .QB(n30917) );
  DFFN img_reg_11__7__6_ ( .D(n12954), .CK(clk), .Q(img[582]), .QB(n30283) );
  DFFN img_reg_11__7__5_ ( .D(n12953), .CK(clk), .Q(img[581]), .QB(n30918) );
  DFFN img_reg_11__6__6_ ( .D(n12942), .CK(clk), .Q(img[590]), .QB(n30439) );
  DFFN img_reg_11__6__5_ ( .D(n12943), .CK(clk), .Q(img[589]), .QB(n30945) );
  DFFN img_reg_11__6__2_ ( .D(n12946), .CK(clk), .Q(img[586]), .QB(n30700) );
  DFFN img_reg_11__5__4_ ( .D(n12936), .CK(clk), .Q(img[596]), .QB(n31899) );
  DFFN img_reg_11__4__6_ ( .D(n12926), .CK(clk), .Q(img[606]), .QB(n30454) );
  DFFN img_reg_11__4__5_ ( .D(n12927), .CK(clk), .Q(img[605]), .QB(n30996) );
  DFFN img_reg_11__4__0_ ( .D(n12932), .CK(clk), .Q(img[600]), .QB(n31668) );
  DFFN img_reg_11__3__5_ ( .D(n12921), .CK(clk), .Q(img[613]), .QB(n30775) );
  DFFN img_reg_11__2__5_ ( .D(n12911), .CK(clk), .Q(img[621]), .QB(n30832) );
  DFFN img_reg_11__1__5_ ( .D(n12905), .CK(clk), .Q(img[629]), .QB(n30972) );
  DFFN img_reg_11__1__3_ ( .D(n12903), .CK(clk), .Q(img[627]), .QB(n31389) );
  DFFN img_reg_11__1__1_ ( .D(n12901), .CK(clk), .Q(img[625]), .QB(n31188) );
  DFFN img_reg_11__1__0_ ( .D(n12908), .CK(clk), .Q(img[624]), .QB(n31636) );
  DFFN img_reg_11__0__5_ ( .D(n12895), .CK(clk), .Q(img[637]), .QB(n30987) );
  DFFN img_reg_11__0__2_ ( .D(n12898), .CK(clk), .Q(img[634]), .QB(n30650) );
  DFFN img_reg_11__9__6_ ( .D(n12970), .CK(clk), .Q(img[566]), .QB(n30438) );
  DFFN img_reg_11__9__5_ ( .D(n12969), .CK(clk), .Q(img[565]), .QB(n30944) );
  DFFN img_reg_13__14__5_ ( .D(n13263), .CK(clk), .Q(img[269]), .QB(n30977) );
  DFFN img_reg_13__14__3_ ( .D(n13265), .CK(clk), .Q(img[267]), .QB(n31406) );
  DFFN img_reg_13__14__0_ ( .D(n13268), .CK(clk), .Q(img[264]), .QB(n31653) );
  DFFN img_reg_12__14__5_ ( .D(n13137), .CK(clk), .Q(img[397]), .QB(n30967) );
  DFFN img_reg_4__14__5_ ( .D(n12113), .CK(clk), .Q(img[1421]), .QB(n30961) );
  DFFN img_reg_4__14__3_ ( .D(n12111), .CK(clk), .Q(img[1419]), .QB(n31411) );
  DFFN img_reg_1__10__1_ ( .D(n11699), .CK(clk), .Q(img[1833]), .QB(n31152) );
  DFFN img_reg_5__11__6_ ( .D(n12218), .CK(clk), .Q(img[1318]), .QB(n30415) );
  DFFN img_reg_2__9__1_ ( .D(n11819), .CK(clk), .Q(img[1713]), .QB(n31154) );
  DFFN img_reg_4__12__6_ ( .D(n12098), .CK(clk), .Q(img[1438]), .QB(n30430) );
  DFFN img_reg_6__11__6_ ( .D(n12342), .CK(clk), .Q(img[1190]), .QB(n30411) );
  DFFN img_reg_1__13__1_ ( .D(n11717), .CK(clk), .Q(img[1809]), .QB(n31150) );
  DFFN img_reg_7__10__3_ ( .D(n12465), .CK(clk), .Q(img[1067]), .QB(n31305) );
  DFFN img_reg_2__9__3_ ( .D(n11817), .CK(clk), .Q(img[1715]), .QB(n31290) );
  DFFN img_reg_3__10__3_ ( .D(n11953), .CK(clk), .Q(img[1579]), .QB(n31301) );
  DFFN img_reg_1__10__3_ ( .D(n11697), .CK(clk), .Q(img[1835]), .QB(n31287) );
  DFFN img_reg_4__12__3_ ( .D(n12095), .CK(clk), .Q(img[1435]), .QB(n31456) );
  DFFN img_reg_14__15__3_ ( .D(n13401), .CK(clk), .Q(img[131]), .QB(n31474) );
  DFFN img_reg_11__10__3_ ( .D(n12977), .CK(clk), .Q(img[555]), .QB(n31317) );
  DFFN img_reg_11__8__3_ ( .D(n12961), .CK(clk), .Q(img[571]), .QB(n31332) );
  DFFN img_reg_11__7__3_ ( .D(n12951), .CK(clk), .Q(img[579]), .QB(n31333) );
  DFFN img_reg_11__6__3_ ( .D(n12945), .CK(clk), .Q(img[587]), .QB(n31434) );
  DFFN img_reg_11__5__3_ ( .D(n12935), .CK(clk), .Q(img[595]), .QB(n31316) );
  DFFN img_reg_11__4__3_ ( .D(n12929), .CK(clk), .Q(img[603]), .QB(n31441) );
  DFFN img_reg_11__3__3_ ( .D(n12919), .CK(clk), .Q(img[611]), .QB(n31482) );
  DFFN img_reg_11__2__3_ ( .D(n12913), .CK(clk), .Q(img[619]), .QB(n31258) );
  DFFN img_reg_11__0__3_ ( .D(n12897), .CK(clk), .Q(img[635]), .QB(n31469) );
  DFFN img_reg_6__11__3_ ( .D(n12345), .CK(clk), .Q(img[1187]), .QB(n31446) );
  DFFN img_reg_3__13__3_ ( .D(n11975), .CK(clk), .Q(img[1555]), .QB(n31304) );
  DFFN img_reg_0__13__3_ ( .D(n11593), .CK(clk), .Q(img[1939]), .QB(n31315) );
  DFFN img_reg_11__9__3_ ( .D(n12967), .CK(clk), .Q(img[563]), .QB(n31433) );
  DFFN img_reg_7__9__3_ ( .D(n12455), .CK(clk), .Q(img[1075]), .QB(n31415) );
  DFFN img_reg_1__9__3_ ( .D(n11687), .CK(clk), .Q(img[1843]), .QB(n31285) );
  DFFN img_reg_5__12__6_ ( .D(n12222), .CK(clk), .Q(img[1310]), .QB(n30418) );
  DFFN img_reg_14__10__1_ ( .D(n13357), .CK(clk), .Q(img[169]), .QB(n31133) );
  DFFN img_reg_14__5__1_ ( .D(n13323), .CK(clk), .Q(img[209]), .QB(n31134) );
  DFFN img_reg_14__12__6_ ( .D(n13378), .CK(clk), .Q(img[158]), .QB(n30422) );
  DFFN img_reg_12__5__1_ ( .D(n13067), .CK(clk), .Q(img[465]), .QB(n31138) );
  DFFN img_reg_14__3__6_ ( .D(n13302), .CK(clk), .Q(img[230]), .QB(n30421) );
  DFFN img_reg_12__3__6_ ( .D(n13046), .CK(clk), .Q(img[486]), .QB(n30425) );
  DFFN img_reg_14__9__3_ ( .D(n13353), .CK(clk), .Q(img[179]), .QB(n31423) );
  DFFN img_reg_14__11__3_ ( .D(n13369), .CK(clk), .Q(img[163]), .QB(n31454) );
  DFFN img_reg_11__8__7_ ( .D(n12957), .CK(clk), .Q(img[575]), .QB(n30164) );
  DFFN img_reg_11__7__7_ ( .D(n12955), .CK(clk), .Q(img[583]), .QB(n30165) );
  DFFN img_reg_0__14__3_ ( .D(n11599), .CK(clk), .Q(img[1931]), .QB(n31311) );
  DFFN img_reg_5__12__3_ ( .D(n12225), .CK(clk), .Q(img[1307]), .QB(n31448) );
  DFFN img_reg_14__13__3_ ( .D(n13385), .CK(clk), .Q(img[147]), .QB(n31273) );
  DFFN img_reg_14__10__3_ ( .D(n13359), .CK(clk), .Q(img[171]), .QB(n31323) );
  DFFN img_reg_14__8__3_ ( .D(n13343), .CK(clk), .Q(img[187]), .QB(n31346) );
  DFFN img_reg_14__7__3_ ( .D(n13337), .CK(clk), .Q(img[195]), .QB(n31347) );
  DFFN img_reg_14__6__3_ ( .D(n13327), .CK(clk), .Q(img[203]), .QB(n31424) );
  DFFN img_reg_14__5__3_ ( .D(n13321), .CK(clk), .Q(img[211]), .QB(n31322) );
  DFFN img_reg_14__12__3_ ( .D(n13375), .CK(clk), .Q(img[155]), .QB(n31487) );
  DFFN img_reg_12__11__3_ ( .D(n13113), .CK(clk), .Q(img[419]), .QB(n31435) );
  DFFN img_reg_12__8__3_ ( .D(n13088), .CK(clk), .Q(img[443]), .QB(n31350) );
  DFFN img_reg_12__7__3_ ( .D(n13081), .CK(clk), .Q(img[451]), .QB(n31351) );
  DFFN img_reg_14__3__3_ ( .D(n13305), .CK(clk), .Q(img[227]), .QB(n31488) );
  DFFN img_reg_14__0__3_ ( .D(n13278), .CK(clk), .Q(img[251]), .QB(n31475) );
  DFFN img_reg_12__3__3_ ( .D(n13049), .CK(clk), .Q(img[483]), .QB(n31492) );
  DFFN img_reg_12__2__3_ ( .D(n13039), .CK(clk), .Q(img[491]), .QB(n31276) );
  DFFN img_reg_14__4__3_ ( .D(n13311), .CK(clk), .Q(img[219]), .QB(n31455) );
  DFFN img_reg_12__4__3_ ( .D(n13055), .CK(clk), .Q(img[475]), .QB(n31436) );
  DFFN img_reg_1__8__3_ ( .D(n11681), .CK(clk), .Q(img[1851]), .QB(n31364) );
  DFFN img_reg_15__8__3_ ( .D(n13473), .CK(clk), .Q(img[59]), .QB(n31334) );
  DFFN img_reg_15__7__3_ ( .D(n13463), .CK(clk), .Q(img[67]), .QB(n31335) );
  DFFN img_reg_15__5__3_ ( .D(n13447), .CK(clk), .Q(img[83]), .QB(n31318) );
  DFFN img_reg_1__12__3_ ( .D(n11713), .CK(clk), .Q(img[1819]), .QB(n31360) );
  DFFN img_reg_15__0__3_ ( .D(n13409), .CK(clk), .Q(img[123]), .QB(n31471) );
  DFFN img_reg_15__2__3_ ( .D(n13425), .CK(clk), .Q(img[107]), .QB(n31260) );
  DFFN img_reg_6__12__3_ ( .D(n12351), .CK(clk), .Q(img[1179]), .QB(n31444) );
  DFFN img_reg_8__7__3_ ( .D(n12569), .CK(clk), .Q(img[963]), .QB(n31345) );
  DFFN img_reg_8__4__3_ ( .D(n12543), .CK(clk), .Q(img[987]), .QB(n31453) );
  DFFN img_reg_8__0__3_ ( .D(n12511), .CK(clk), .Q(img[1019]), .QB(n31473) );
  DFFN img_reg_14__8__7_ ( .D(n13347), .CK(clk), .Q(img[191]), .QB(n30178) );
  DFFN img_reg_14__7__7_ ( .D(n13333), .CK(clk), .Q(img[199]), .QB(n30179) );
  DFFN img_reg_12__7__7_ ( .D(n13077), .CK(clk), .Q(img[455]), .QB(n30183) );
  DFFN img_reg_6__8__7_ ( .D(n12323), .CK(clk), .Q(img[1215]), .QB(n30170) );
  DFFN img_reg_11__2__4_ ( .D(n12912), .CK(clk), .Q(img[620]), .QB(n31868) );
  DFFN img_reg_5__13__4_ ( .D(n12232), .CK(clk), .Q(img[1300]), .QB(n31877) );
  DFFN img_reg_14__2__4_ ( .D(n13296), .CK(clk), .Q(img[236]), .QB(n31882) );
  DFFN img_reg_14__13__4_ ( .D(n13384), .CK(clk), .Q(img[148]), .QB(n31881) );
  DFFN img_reg_12__2__4_ ( .D(n13040), .CK(clk), .Q(img[492]), .QB(n31886) );
  DFFN img_reg_15__2__4_ ( .D(n13424), .CK(clk), .Q(img[108]), .QB(n31870) );
  DFFN img_reg_6__10__4_ ( .D(n12336), .CK(clk), .Q(img[1196]), .QB(n31871) );
  DFFN img_reg_7__10__2_ ( .D(n12466), .CK(clk), .Q(img[1066]), .QB(n30620) );
  DFFN img_reg_3__10__2_ ( .D(n11954), .CK(clk), .Q(img[1578]), .QB(n30571) );
  DFFN img_reg_5__11__2_ ( .D(n12214), .CK(clk), .Q(img[1314]), .QB(n30722) );
  DFFN img_reg_5__11__0_ ( .D(n12220), .CK(clk), .Q(img[1312]), .QB(n31677) );
  DFFN img_reg_1__10__2_ ( .D(n11698), .CK(clk), .Q(img[1834]), .QB(n30555) );
  DFFN img_reg_1__10__0_ ( .D(n11700), .CK(clk), .Q(img[1832]), .QB(n31604) );
  DFFN img_reg_2__9__2_ ( .D(n11818), .CK(clk), .Q(img[1714]), .QB(n30567) );
  DFFN img_reg_4__12__2_ ( .D(n12094), .CK(clk), .Q(img[1434]), .QB(n30730) );
  DFFN img_reg_4__12__0_ ( .D(n12100), .CK(clk), .Q(img[1432]), .QB(n31687) );
  DFFN img_reg_14__15__0_ ( .D(n13404), .CK(clk), .Q(img[128]), .QB(n31566) );
  DFFN img_reg_11__10__2_ ( .D(n12978), .CK(clk), .Q(img[554]), .QB(n30591) );
  DFFN img_reg_11__10__0_ ( .D(n12980), .CK(clk), .Q(img[552]), .QB(n31989) );
  DFFN img_reg_11__8__2_ ( .D(n12962), .CK(clk), .Q(img[570]), .QB(n31993) );
  DFFN img_reg_11__8__0_ ( .D(n12964), .CK(clk), .Q(img[568]), .QB(n31509) );
  DFFN img_reg_11__7__0_ ( .D(n12956), .CK(clk), .Q(img[576]), .QB(n31510) );
  DFFN img_reg_11__6__0_ ( .D(n12948), .CK(clk), .Q(img[584]), .QB(n31713) );
  DFFN img_reg_11__5__2_ ( .D(n12934), .CK(clk), .Q(img[594]), .QB(n30592) );
  DFFN img_reg_11__5__0_ ( .D(n12940), .CK(clk), .Q(img[592]), .QB(n31700) );
  DFFN img_reg_11__4__2_ ( .D(n12930), .CK(clk), .Q(img[602]), .QB(n30742) );
  DFFN img_reg_11__3__2_ ( .D(n12918), .CK(clk), .Q(img[610]), .QB(n30745) );
  DFFN img_reg_11__3__0_ ( .D(n12924), .CK(clk), .Q(img[608]), .QB(n31728) );
  DFFN img_reg_11__2__2_ ( .D(n12914), .CK(clk), .Q(img[618]), .QB(n30626) );
  DFFN img_reg_11__2__0_ ( .D(n12916), .CK(clk), .Q(img[616]), .QB(n31574) );
  DFFN img_reg_11__1__2_ ( .D(n12902), .CK(clk), .Q(img[626]), .QB(n30528) );
  DFFN img_reg_11__0__0_ ( .D(n12900), .CK(clk), .Q(img[632]), .QB(n31559) );
  DFFN img_reg_6__11__2_ ( .D(n12346), .CK(clk), .Q(img[1186]), .QB(n30718) );
  DFFN img_reg_6__11__0_ ( .D(n12348), .CK(clk), .Q(img[1184]), .QB(n31673) );
  DFFN img_reg_5__13__2_ ( .D(n12230), .CK(clk), .Q(img[1298]), .QB(n30599) );
  DFFN img_reg_3__13__2_ ( .D(n11974), .CK(clk), .Q(img[1554]), .QB(n30573) );
  DFFN img_reg_1__13__2_ ( .D(n11718), .CK(clk), .Q(img[1810]), .QB(n30557) );
  DFFN img_reg_0__13__2_ ( .D(n11594), .CK(clk), .Q(img[1938]), .QB(n30585) );
  DFFN img_reg_11__9__0_ ( .D(n12972), .CK(clk), .Q(img[560]), .QB(n31712) );
  DFFN img_reg_13__14__2_ ( .D(n13266), .CK(clk), .Q(img[266]), .QB(n30545) );
  DFFN img_reg_12__14__2_ ( .D(n13134), .CK(clk), .Q(img[394]), .QB(n30547) );
  DFFN img_reg_4__14__0_ ( .D(n12116), .CK(clk), .Q(img[1416]), .QB(n31659) );
  DFFN img_reg_7__9__2_ ( .D(n12454), .CK(clk), .Q(img[1074]), .QB(n30579) );
  DFFN img_reg_5__9__2_ ( .D(n12198), .CK(clk), .Q(img[1330]), .QB(n30536) );
  DFFN img_reg_1__9__0_ ( .D(n11692), .CK(clk), .Q(img[1840]), .QB(n31600) );
  DFFN img_reg_14__9__2_ ( .D(n13354), .CK(clk), .Q(img[178]), .QB(n30705) );
  DFFN img_reg_14__11__2_ ( .D(n13370), .CK(clk), .Q(img[162]), .QB(n30724) );
  DFFN img_reg_14__9__0_ ( .D(n13356), .CK(clk), .Q(img[176]), .QB(n31718) );
  DFFN img_reg_14__2__2_ ( .D(n13294), .CK(clk), .Q(img[234]), .QB(n30632) );
  DFFN img_reg_14__11__0_ ( .D(n13372), .CK(clk), .Q(img[160]), .QB(n31681) );
  DFFN img_reg_0__14__2_ ( .D(n11598), .CK(clk), .Q(img[1930]), .QB(n30590) );
  DFFN img_reg_5__12__2_ ( .D(n12226), .CK(clk), .Q(img[1306]), .QB(n30720) );
  DFFN img_reg_5__12__0_ ( .D(n12228), .CK(clk), .Q(img[1304]), .QB(n31675) );
  DFFN img_reg_0__12__2_ ( .D(n11582), .CK(clk), .Q(img[1946]), .QB(n30643) );
  DFFN img_reg_0__12__0_ ( .D(n11588), .CK(clk), .Q(img[1944]), .QB(n31553) );
  DFFN img_reg_14__13__2_ ( .D(n13386), .CK(clk), .Q(img[146]), .QB(n30633) );
  DFFN img_reg_14__13__0_ ( .D(n13388), .CK(clk), .Q(img[144]), .QB(n31587) );
  DFFN img_reg_14__10__2_ ( .D(n13358), .CK(clk), .Q(img[170]), .QB(n30605) );
  DFFN img_reg_14__10__0_ ( .D(n13364), .CK(clk), .Q(img[168]), .QB(n31698) );
  DFFN img_reg_14__8__2_ ( .D(n13342), .CK(clk), .Q(img[186]), .QB(n30766) );
  DFFN img_reg_14__8__0_ ( .D(n13348), .CK(clk), .Q(img[184]), .QB(n31523) );
  DFFN img_reg_14__7__2_ ( .D(n13338), .CK(clk), .Q(img[194]), .QB(n30767) );
  DFFN img_reg_14__7__0_ ( .D(n13340), .CK(clk), .Q(img[192]), .QB(n31524) );
  DFFN img_reg_14__6__0_ ( .D(n13332), .CK(clk), .Q(img[200]), .QB(n31719) );
  DFFN img_reg_14__5__2_ ( .D(n13322), .CK(clk), .Q(img[210]), .QB(n30606) );
  DFFN img_reg_14__5__0_ ( .D(n13324), .CK(clk), .Q(img[208]), .QB(n31699) );
  DFFN img_reg_14__12__2_ ( .D(n13374), .CK(clk), .Q(img[154]), .QB(n30752) );
  DFFN img_reg_14__12__0_ ( .D(n13380), .CK(clk), .Q(img[152]), .QB(n31733) );
  DFFN img_reg_12__11__0_ ( .D(n13116), .CK(clk), .Q(img[416]), .QB(n31685) );
  DFFN img_reg_12__10__2_ ( .D(n13102), .CK(clk), .Q(img[426]), .QB(n30609) );
  DFFN img_reg_12__7__2_ ( .D(n13082), .CK(clk), .Q(img[450]), .QB(n30771) );
  DFFN img_reg_12__7__0_ ( .D(n13084), .CK(clk), .Q(img[448]), .QB(n31528) );
  DFFN img_reg_12__5__2_ ( .D(n13066), .CK(clk), .Q(img[466]), .QB(n30610) );
  DFFN img_reg_12__5__0_ ( .D(n13068), .CK(clk), .Q(img[464]), .QB(n31708) );
  DFFN img_reg_14__3__2_ ( .D(n13306), .CK(clk), .Q(img[226]), .QB(n30751) );
  DFFN img_reg_14__3__0_ ( .D(n13308), .CK(clk), .Q(img[224]), .QB(n31734) );
  DFFN img_reg_14__1__2_ ( .D(n13290), .CK(clk), .Q(img[242]), .QB(n30542) );
  DFFN img_reg_12__3__2_ ( .D(n13050), .CK(clk), .Q(img[482]), .QB(n30755) );
  DFFN img_reg_12__3__0_ ( .D(n13052), .CK(clk), .Q(img[480]), .QB(n31738) );
  DFFN img_reg_12__2__2_ ( .D(n13038), .CK(clk), .Q(img[490]), .QB(n30634) );
  DFFN img_reg_12__2__0_ ( .D(n13044), .CK(clk), .Q(img[488]), .QB(n31592) );
  DFFN img_reg_12__1__2_ ( .D(n13034), .CK(clk), .Q(img[498]), .QB(n30546) );
  DFFN img_reg_14__4__2_ ( .D(n13310), .CK(clk), .Q(img[218]), .QB(n30725) );
  DFFN img_reg_14__4__0_ ( .D(n13316), .CK(clk), .Q(img[216]), .QB(n31682) );
  DFFN img_reg_12__4__2_ ( .D(n13054), .CK(clk), .Q(img[474]), .QB(n30729) );
  DFFN img_reg_12__4__0_ ( .D(n13060), .CK(clk), .Q(img[472]), .QB(n31686) );
  DFFN img_reg_1__8__0_ ( .D(n11684), .CK(clk), .Q(img[1848]), .QB(n31507) );
  DFFN img_reg_0__8__2_ ( .D(n11550), .CK(clk), .Q(img[1978]), .QB(n30645) );
  DFFN img_reg_0__8__0_ ( .D(n11556), .CK(clk), .Q(img[1976]), .QB(n31557) );
  DFFN img_reg_3__12__0_ ( .D(n11972), .CK(clk), .Q(img[1560]), .QB(n31541) );
  DFFN img_reg_15__4__0_ ( .D(n13444), .CK(clk), .Q(img[88]), .QB(n31670) );
  DFFN img_reg_6__8__0_ ( .D(n12324), .CK(clk), .Q(img[1208]), .QB(n31499) );
  DFFN img_reg_12__0__3_ ( .D(n13023), .CK(clk), .Q(img[507]), .QB(n31467) );
  DFFN img_reg_3__10__6_ ( .D(n11950), .CK(clk), .Q(img[1582]), .QB(n30387) );
  DFFN img_reg_3__10__1_ ( .D(n11955), .CK(clk), .Q(img[1577]), .QB(n31168) );
  DFFN img_reg_2__9__6_ ( .D(n11814), .CK(clk), .Q(img[1718]), .QB(n30383) );
  DFFN img_reg_1__10__6_ ( .D(n11694), .CK(clk), .Q(img[1838]), .QB(n30371) );
  DFFN img_reg_7__10__6_ ( .D(n12462), .CK(clk), .Q(img[1070]), .QB(n30493) );
  DFFN img_reg_5__11__1_ ( .D(n12213), .CK(clk), .Q(img[1313]), .QB(n31084) );
  DFFN img_reg_4__12__1_ ( .D(n12093), .CK(clk), .Q(img[1433]), .QB(n31093) );
  DFFN img_reg_14__15__6_ ( .D(n13398), .CK(clk), .Q(img[134]), .QB(n30477) );
  DFFN img_reg_14__15__1_ ( .D(n13403), .CK(clk), .Q(img[129]), .QB(n31026) );
  DFFN img_reg_11__10__6_ ( .D(n12974), .CK(clk), .Q(img[558]), .QB(n30495) );
  DFFN img_reg_11__10__1_ ( .D(n12979), .CK(clk), .Q(img[553]), .QB(n31119) );
  DFFN img_reg_11__8__6_ ( .D(n12958), .CK(clk), .Q(img[574]), .QB(n31994) );
  DFFN img_reg_11__7__1_ ( .D(n12949), .CK(clk), .Q(img[577]), .QB(n31229) );
  DFFN img_reg_11__6__1_ ( .D(n12947), .CK(clk), .Q(img[585]), .QB(n31214) );
  DFFN img_reg_11__5__6_ ( .D(n12938), .CK(clk), .Q(img[598]), .QB(n30494) );
  DFFN img_reg_11__5__1_ ( .D(n12933), .CK(clk), .Q(img[593]), .QB(n31120) );
  DFFN img_reg_11__4__1_ ( .D(n12931), .CK(clk), .Q(img[601]), .QB(n31991) );
  DFFN img_reg_11__3__6_ ( .D(n12922), .CK(clk), .Q(img[614]), .QB(n30407) );
  DFFN img_reg_11__3__1_ ( .D(n12917), .CK(clk), .Q(img[609]), .QB(n31104) );
  DFFN img_reg_11__2__6_ ( .D(n12910), .CK(clk), .Q(img[622]), .QB(n30514) );
  DFFN img_reg_11__2__1_ ( .D(n12915), .CK(clk), .Q(img[617]), .QB(n31243) );
  DFFN img_reg_11__1__6_ ( .D(n12906), .CK(clk), .Q(img[630]), .QB(n30345) );
  DFFN img_reg_11__0__6_ ( .D(n12894), .CK(clk), .Q(img[638]), .QB(n30472) );
  DFFN img_reg_11__0__1_ ( .D(n12899), .CK(clk), .Q(img[633]), .QB(n31011) );
  DFFN img_reg_6__11__1_ ( .D(n12347), .CK(clk), .Q(img[1185]), .QB(n31080) );
  DFFN img_reg_5__13__6_ ( .D(n12234), .CK(clk), .Q(img[1302]), .QB(n30482) );
  DFFN img_reg_3__13__6_ ( .D(n11978), .CK(clk), .Q(img[1558]), .QB(n30389) );
  DFFN img_reg_1__13__6_ ( .D(n11722), .CK(clk), .Q(img[1814]), .QB(n30373) );
  DFFN img_reg_0__13__6_ ( .D(n11590), .CK(clk), .Q(img[1942]), .QB(n30401) );
  DFFN img_reg_11__9__1_ ( .D(n12965), .CK(clk), .Q(img[561]), .QB(n31213) );
  DFFN img_reg_13__14__6_ ( .D(n13262), .CK(clk), .Q(img[270]), .QB(n30360) );
  DFFN img_reg_13__14__1_ ( .D(n13267), .CK(clk), .Q(img[265]), .QB(n31197) );
  DFFN img_reg_12__14__6_ ( .D(n13138), .CK(clk), .Q(img[398]), .QB(n30362) );
  DFFN img_reg_12__14__1_ ( .D(n13133), .CK(clk), .Q(img[393]), .QB(n31199) );
  DFFN img_reg_4__14__6_ ( .D(n12114), .CK(clk), .Q(img[1422]), .QB(n30366) );
  DFFN img_reg_4__14__1_ ( .D(n12109), .CK(clk), .Q(img[1417]), .QB(n31203) );
  DFFN img_reg_5__9__6_ ( .D(n12202), .CK(clk), .Q(img[1334]), .QB(n30352) );
  DFFN img_reg_5__9__1_ ( .D(n12197), .CK(clk), .Q(img[1329]), .QB(n31191) );
  DFFN img_reg_14__11__6_ ( .D(n13366), .CK(clk), .Q(img[166]), .QB(n30459) );
  DFFN img_reg_14__11__1_ ( .D(n13371), .CK(clk), .Q(img[161]), .QB(n31088) );
  DFFN img_reg_14__9__1_ ( .D(n13355), .CK(clk), .Q(img[177]), .QB(n31219) );
  DFFN img_reg_14__2__6_ ( .D(n13298), .CK(clk), .Q(img[238]), .QB(n30520) );
  DFFN img_reg_14__2__1_ ( .D(n13293), .CK(clk), .Q(img[233]), .QB(n31249) );
  DFFN img_reg_0__14__6_ ( .D(n11602), .CK(clk), .Q(img[1934]), .QB(n30405) );
  DFFN img_reg_5__12__1_ ( .D(n12227), .CK(clk), .Q(img[1305]), .QB(n31081) );
  DFFN img_reg_0__12__6_ ( .D(n11586), .CK(clk), .Q(img[1950]), .QB(n30338) );
  DFFN img_reg_0__12__1_ ( .D(n11581), .CK(clk), .Q(img[1945]), .QB(n31068) );
  DFFN img_reg_14__13__1_ ( .D(n13387), .CK(clk), .Q(img[145]), .QB(n31250) );
  DFFN img_reg_14__10__6_ ( .D(n13362), .CK(clk), .Q(img[174]), .QB(n30505) );
  DFFN img_reg_14__8__6_ ( .D(n13346), .CK(clk), .Q(img[190]), .QB(n30296) );
  DFFN img_reg_14__8__1_ ( .D(n13341), .CK(clk), .Q(img[185]), .QB(n31236) );
  DFFN img_reg_14__7__6_ ( .D(n13334), .CK(clk), .Q(img[198]), .QB(n30297) );
  DFFN img_reg_14__7__1_ ( .D(n13339), .CK(clk), .Q(img[193]), .QB(n31235) );
  DFFN img_reg_14__6__6_ ( .D(n13330), .CK(clk), .Q(img[206]), .QB(n30445) );
  DFFN img_reg_14__5__6_ ( .D(n13318), .CK(clk), .Q(img[214]), .QB(n30504) );
  DFFN img_reg_14__12__1_ ( .D(n13373), .CK(clk), .Q(img[153]), .QB(n31111) );
  DFFN img_reg_12__11__6_ ( .D(n13110), .CK(clk), .Q(img[422]), .QB(n30463) );
  DFFN img_reg_12__11__1_ ( .D(n13115), .CK(clk), .Q(img[417]), .QB(n31092) );
  DFFN img_reg_12__10__6_ ( .D(n13106), .CK(clk), .Q(img[430]), .QB(n30509) );
  DFFN img_reg_12__7__6_ ( .D(n13078), .CK(clk), .Q(img[454]), .QB(n30301) );
  DFFN img_reg_12__7__1_ ( .D(n13083), .CK(clk), .Q(img[449]), .QB(n31239) );
  DFFN img_reg_12__5__6_ ( .D(n13062), .CK(clk), .Q(img[470]), .QB(n30508) );
  DFFN img_reg_14__3__1_ ( .D(n13307), .CK(clk), .Q(img[225]), .QB(n31110) );
  DFFN img_reg_14__1__6_ ( .D(n13286), .CK(clk), .Q(img[246]), .QB(n30359) );
  DFFN img_reg_14__1__1_ ( .D(n13291), .CK(clk), .Q(img[241]), .QB(n31196) );
  DFFN img_reg_14__0__6_ ( .D(n13281), .CK(clk), .Q(img[254]), .QB(n30478) );
  DFFN img_reg_14__0__1_ ( .D(n13283), .CK(clk), .Q(img[249]), .QB(n31025) );
  DFFN img_reg_12__3__1_ ( .D(n13051), .CK(clk), .Q(img[481]), .QB(n31114) );
  DFFN img_reg_12__2__1_ ( .D(n13037), .CK(clk), .Q(img[489]), .QB(n31253) );
  DFFN img_reg_12__1__6_ ( .D(n13030), .CK(clk), .Q(img[502]), .QB(n30363) );
  DFFN img_reg_12__1__1_ ( .D(n13035), .CK(clk), .Q(img[497]), .QB(n31200) );
  DFFN img_reg_14__4__6_ ( .D(n13314), .CK(clk), .Q(img[222]), .QB(n30460) );
  DFFN img_reg_14__4__1_ ( .D(n13309), .CK(clk), .Q(img[217]), .QB(n31087) );
  DFFN img_reg_12__4__6_ ( .D(n13058), .CK(clk), .Q(img[478]), .QB(n30464) );
  DFFN img_reg_12__4__1_ ( .D(n13053), .CK(clk), .Q(img[473]), .QB(n31091) );
  DFFN img_reg_1__8__6_ ( .D(n11678), .CK(clk), .Q(img[1854]), .QB(n30314) );
  DFFN img_reg_1__8__1_ ( .D(n11683), .CK(clk), .Q(img[1849]), .QB(n31042) );
  DFFN img_reg_0__8__6_ ( .D(n11554), .CK(clk), .Q(img[1982]), .QB(n30342) );
  DFFN img_reg_0__8__1_ ( .D(n11549), .CK(clk), .Q(img[1977]), .QB(n31070) );
  DFFN img_reg_6__8__6_ ( .D(n12322), .CK(clk), .Q(img[1214]), .QB(n30288) );
  DFFN img_reg_6__8__1_ ( .D(n12317), .CK(clk), .Q(img[1209]), .QB(n31015) );
  DFFN img_reg_7__10__7_ ( .D(n12461), .CK(clk), .Q(img[1071]), .QB(n30221) );
  DFFN img_reg_1__10__7_ ( .D(n11693), .CK(clk), .Q(img[1839]), .QB(n30065) );
  DFFN img_reg_5__11__7_ ( .D(n12219), .CK(clk), .Q(img[1319]), .QB(n30109) );
  DFFN img_reg_2__9__7_ ( .D(n11813), .CK(clk), .Q(img[1719]), .QB(n30079) );
  DFFN img_reg_4__12__7_ ( .D(n12099), .CK(clk), .Q(img[1439]), .QB(n30124) );
  DFFN img_reg_14__15__7_ ( .D(n13397), .CK(clk), .Q(img[135]), .QB(n30274) );
  DFFN img_reg_11__10__7_ ( .D(n12973), .CK(clk), .Q(img[559]), .QB(n30226) );
  DFFN img_reg_11__6__7_ ( .D(n12941), .CK(clk), .Q(img[591]), .QB(n30038) );
  DFFN img_reg_11__5__7_ ( .D(n12939), .CK(clk), .Q(img[599]), .QB(n30225) );
  DFFN img_reg_11__4__7_ ( .D(n12925), .CK(clk), .Q(img[607]), .QB(n30243) );
  DFFN img_reg_11__3__7_ ( .D(n12923), .CK(clk), .Q(img[615]), .QB(n30101) );
  DFFN img_reg_11__2__7_ ( .D(n12909), .CK(clk), .Q(img[623]), .QB(n30194) );
  DFFN img_reg_11__1__7_ ( .D(n12907), .CK(clk), .Q(img[631]), .QB(n30256) );
  DFFN img_reg_11__0__7_ ( .D(n12893), .CK(clk), .Q(img[639]), .QB(n30269) );
  DFFN img_reg_6__11__7_ ( .D(n12341), .CK(clk), .Q(img[1191]), .QB(n30105) );
  DFFN img_reg_3__13__7_ ( .D(n11979), .CK(clk), .Q(img[1559]), .QB(n30083) );
  DFFN img_reg_1__13__7_ ( .D(n11723), .CK(clk), .Q(img[1815]), .QB(n30067) );
  DFFN img_reg_0__13__7_ ( .D(n11589), .CK(clk), .Q(img[1943]), .QB(n30095) );
  DFFN img_reg_11__9__7_ ( .D(n12971), .CK(clk), .Q(img[567]), .QB(n30037) );
  DFFN img_reg_13__14__7_ ( .D(n13261), .CK(clk), .Q(img[271]), .QB(n30261) );
  DFFN img_reg_4__14__7_ ( .D(n12115), .CK(clk), .Q(img[1423]), .QB(n30058) );
  DFFN img_reg_5__9__7_ ( .D(n12203), .CK(clk), .Q(img[1335]), .QB(n30048) );
  DFFN img_reg_14__9__7_ ( .D(n13349), .CK(clk), .Q(img[183]), .QB(n30052) );
  DFFN img_reg_14__11__7_ ( .D(n13365), .CK(clk), .Q(img[167]), .QB(n30248) );
  DFFN img_reg_14__2__7_ ( .D(n13299), .CK(clk), .Q(img[239]), .QB(n30208) );
  DFFN img_reg_0__14__7_ ( .D(n11603), .CK(clk), .Q(img[1935]), .QB(n30097) );
  DFFN img_reg_5__12__7_ ( .D(n12221), .CK(clk), .Q(img[1311]), .QB(n30112) );
  DFFN img_reg_2__12__7_ ( .D(n11843), .CK(clk), .Q(img[1695]), .QB(n30143) );
  DFFN img_reg_0__12__7_ ( .D(n11587), .CK(clk), .Q(img[1951]), .QB(n30163) );
  DFFN img_reg_14__6__7_ ( .D(n13331), .CK(clk), .Q(img[207]), .QB(n30053) );
  DFFN img_reg_14__5__7_ ( .D(n13317), .CK(clk), .Q(img[215]), .QB(n30229) );
  DFFN img_reg_14__12__7_ ( .D(n13379), .CK(clk), .Q(img[159]), .QB(n30116) );
  DFFN img_reg_12__11__7_ ( .D(n13109), .CK(clk), .Q(img[423]), .QB(n30250) );
  DFFN img_reg_12__10__7_ ( .D(n13107), .CK(clk), .Q(img[431]), .QB(n30234) );
  DFFN img_reg_12__5__7_ ( .D(n13061), .CK(clk), .Q(img[471]), .QB(n30233) );
  DFFN img_reg_14__3__7_ ( .D(n13301), .CK(clk), .Q(img[231]), .QB(n30115) );
  DFFN img_reg_14__1__7_ ( .D(n13285), .CK(clk), .Q(img[247]), .QB(n30260) );
  DFFN img_reg_14__0__7_ ( .D(n13282), .CK(clk), .Q(img[255]), .QB(n30275) );
  DFFN img_reg_12__3__7_ ( .D(n13045), .CK(clk), .Q(img[487]), .QB(n30119) );
  DFFN img_reg_12__1__7_ ( .D(n13029), .CK(clk), .Q(img[503]), .QB(n30264) );
  DFFN img_reg_14__4__7_ ( .D(n13315), .CK(clk), .Q(img[223]), .QB(n30249) );
  DFFN img_reg_12__4__7_ ( .D(n13059), .CK(clk), .Q(img[479]), .QB(n30251) );
  DFFN img_reg_1__8__7_ ( .D(n11677), .CK(clk), .Q(img[1855]), .QB(n30128) );
  DFFN img_reg_15__11__7_ ( .D(n13499), .CK(clk), .Q(img[39]), .QB(n30244) );
  DFFN img_reg_12__12__7_ ( .D(n13123), .CK(clk), .Q(img[415]), .QB(n30120) );
  DFFN img_reg_3__12__7_ ( .D(n11965), .CK(clk), .Q(img[1567]), .QB(n30151) );
  DFFN img_reg_1__12__7_ ( .D(n11709), .CK(clk), .Q(img[1823]), .QB(n30135) );
  DFFN img_reg_15__4__7_ ( .D(n13437), .CK(clk), .Q(img[95]), .QB(n30245) );
  DFFN img_reg_10__12__7_ ( .D(n12867), .CK(clk), .Q(img[671]), .QB(n30127) );
  DFFN img_reg_9__12__7_ ( .D(n12733), .CK(clk), .Q(img[799]), .QB(n30125) );
  DFFN img_reg_8__4__7_ ( .D(n12547), .CK(clk), .Q(img[991]), .QB(n30247) );
  DFFN img_reg_8__1__7_ ( .D(n12517), .CK(clk), .Q(img[1015]), .QB(n30258) );
  DFFN img_reg_7__10__4_ ( .D(n12464), .CK(clk), .Q(img[1068]), .QB(n31894) );
  DFFN img_reg_2__9__4_ ( .D(n11816), .CK(clk), .Q(img[1716]), .QB(n31783) );
  DFFN img_reg_5__11__4_ ( .D(n12216), .CK(clk), .Q(img[1316]), .QB(n31929) );
  DFFN img_reg_3__10__4_ ( .D(n11952), .CK(clk), .Q(img[1580]), .QB(n31785) );
  DFFN img_reg_1__10__4_ ( .D(n11696), .CK(clk), .Q(img[1836]), .QB(n31769) );
  DFFN img_reg_14__15__4_ ( .D(n13400), .CK(clk), .Q(img[132]), .QB(n31980) );
  DFFN img_reg_11__10__4_ ( .D(n12976), .CK(clk), .Q(img[556]), .QB(n31898) );
  DFFN img_reg_11__8__4_ ( .D(n12960), .CK(clk), .Q(img[572]), .QB(n31806) );
  DFFN img_reg_11__7__4_ ( .D(n12952), .CK(clk), .Q(img[580]), .QB(n31805) );
  DFFN img_reg_11__6__4_ ( .D(n12944), .CK(clk), .Q(img[588]), .QB(n31743) );
  DFFN img_reg_11__4__4_ ( .D(n12928), .CK(clk), .Q(img[604]), .QB(n31988) );
  DFFN img_reg_11__3__4_ ( .D(n12920), .CK(clk), .Q(img[612]), .QB(n31944) );
  DFFN img_reg_11__1__4_ ( .D(n12904), .CK(clk), .Q(img[628]), .QB(n31946) );
  DFFN img_reg_11__0__4_ ( .D(n12896), .CK(clk), .Q(img[636]), .QB(n31975) );
  DFFN img_reg_6__11__4_ ( .D(n12344), .CK(clk), .Q(img[1188]), .QB(n31921) );
  DFFN img_reg_7__13__4_ ( .D(n12487), .CK(clk), .Q(img[1044]), .QB(n31896) );
  DFFN img_reg_3__13__4_ ( .D(n11976), .CK(clk), .Q(img[1556]), .QB(n31787) );
  DFFN img_reg_2__13__4_ ( .D(n11848), .CK(clk), .Q(img[1684]), .QB(n31779) );
  DFFN img_reg_1__13__4_ ( .D(n11720), .CK(clk), .Q(img[1812]), .QB(n31771) );
  DFFN img_reg_11__9__4_ ( .D(n12968), .CK(clk), .Q(img[564]), .QB(n31742) );
  DFFN img_reg_13__14__4_ ( .D(n13264), .CK(clk), .Q(img[268]), .QB(n31953) );
  DFFN img_reg_12__14__4_ ( .D(n13136), .CK(clk), .Q(img[396]), .QB(n31955) );
  DFFN img_reg_4__14__4_ ( .D(n12112), .CK(clk), .Q(img[1420]), .QB(n31762) );
  DFFN img_reg_7__9__4_ ( .D(n12456), .CK(clk), .Q(img[1076]), .QB(n31795) );
  DFFN img_reg_5__9__4_ ( .D(n12200), .CK(clk), .Q(img[1332]), .QB(n31752) );
  DFFN img_reg_1__9__4_ ( .D(n11688), .CK(clk), .Q(img[1844]), .QB(n31775) );
  DFFN img_reg_14__11__4_ ( .D(n13368), .CK(clk), .Q(img[164]), .QB(n31966) );
  DFFN img_reg_14__9__4_ ( .D(n13352), .CK(clk), .Q(img[180]), .QB(n31756) );
  DFFN img_reg_7__14__4_ ( .D(n12496), .CK(clk), .Q(img[1036]), .QB(n31793) );
  DFFN img_reg_2__14__4_ ( .D(n11856), .CK(clk), .Q(img[1676]), .QB(n31781) );
  DFFN img_reg_0__14__4_ ( .D(n11600), .CK(clk), .Q(img[1932]), .QB(n31801) );
  DFFN img_reg_5__12__4_ ( .D(n12224), .CK(clk), .Q(img[1308]), .QB(n31931) );
  DFFN img_reg_2__12__4_ ( .D(n11840), .CK(clk), .Q(img[1692]), .QB(n31841) );
  DFFN img_reg_14__8__4_ ( .D(n13344), .CK(clk), .Q(img[188]), .QB(n31820) );
  DFFN img_reg_14__7__4_ ( .D(n13336), .CK(clk), .Q(img[196]), .QB(n31819) );
  DFFN img_reg_14__6__4_ ( .D(n13328), .CK(clk), .Q(img[204]), .QB(n31757) );
  DFFN img_reg_14__12__4_ ( .D(n13376), .CK(clk), .Q(img[156]), .QB(n31937) );
  DFFN img_reg_12__11__4_ ( .D(n13112), .CK(clk), .Q(img[420]), .QB(n31970) );
  DFFN img_reg_12__8__4_ ( .D(n13089), .CK(clk), .Q(img[444]), .QB(n31824) );
  DFFN img_reg_12__7__4_ ( .D(n13080), .CK(clk), .Q(img[452]), .QB(n31823) );
  DFFN img_reg_12__5__4_ ( .D(n13064), .CK(clk), .Q(img[468]), .QB(n31909) );
  DFFN img_reg_14__3__4_ ( .D(n13304), .CK(clk), .Q(img[228]), .QB(n31938) );
  DFFN img_reg_14__1__4_ ( .D(n13288), .CK(clk), .Q(img[244]), .QB(n31952) );
  DFFN img_reg_14__0__4_ ( .D(n13279), .CK(clk), .Q(img[252]), .QB(n31981) );
  DFFN img_reg_12__3__4_ ( .D(n13048), .CK(clk), .Q(img[484]), .QB(n31940) );
  DFFN img_reg_12__1__4_ ( .D(n13032), .CK(clk), .Q(img[500]), .QB(n31956) );
  DFFN img_reg_14__4__4_ ( .D(n13312), .CK(clk), .Q(img[220]), .QB(n31965) );
  DFFN img_reg_1__8__4_ ( .D(n11680), .CK(clk), .Q(img[1852]), .QB(n31838) );
  DFFN img_reg_0__8__4_ ( .D(n11552), .CK(clk), .Q(img[1980]), .QB(n31866) );
  DFFN img_reg_15__12__4_ ( .D(n13504), .CK(clk), .Q(img[28]), .QB(n31941) );
  DFFN img_reg_15__11__4_ ( .D(n13496), .CK(clk), .Q(img[36]), .QB(n31962) );
  DFFN img_reg_15__8__4_ ( .D(n13472), .CK(clk), .Q(img[60]), .QB(n31808) );
  DFFN img_reg_15__7__4_ ( .D(n13464), .CK(clk), .Q(img[68]), .QB(n31807) );
  DFFN img_reg_15__6__4_ ( .D(n13456), .CK(clk), .Q(img[76]), .QB(n31745) );
  DFFN img_reg_12__12__4_ ( .D(n13120), .CK(clk), .Q(img[412]), .QB(n31939) );
  DFFN img_reg_7__12__4_ ( .D(n12480), .CK(clk), .Q(img[1052]), .QB(n31917) );
  DFFN img_reg_3__12__4_ ( .D(n11968), .CK(clk), .Q(img[1564]), .QB(n31849) );
  DFFN img_reg_1__12__4_ ( .D(n11712), .CK(clk), .Q(img[1820]), .QB(n31833) );
  DFFN img_reg_15__4__4_ ( .D(n13440), .CK(clk), .Q(img[92]), .QB(n31961) );
  DFFN img_reg_15__3__4_ ( .D(n13432), .CK(clk), .Q(img[100]), .QB(n31942) );
  DFFN img_reg_15__1__4_ ( .D(n13416), .CK(clk), .Q(img[116]), .QB(n31948) );
  DFFN img_reg_11__12__4_ ( .D(n12992), .CK(clk), .Q(img[540]), .QB(n31943) );
  DFFN img_reg_10__12__4_ ( .D(n12864), .CK(clk), .Q(img[668]), .QB(n31919) );
  DFFN img_reg_9__12__4_ ( .D(n12736), .CK(clk), .Q(img[796]), .QB(n31927) );
  DFFN img_reg_8__12__4_ ( .D(n12608), .CK(clk), .Q(img[924]), .QB(n31925) );
  DFFN img_reg_6__12__4_ ( .D(n12352), .CK(clk), .Q(img[1180]), .QB(n31923) );
  DFFN img_reg_6__8__4_ ( .D(n12320), .CK(clk), .Q(img[1212]), .QB(n31812) );
  DFFN img_reg_8__7__4_ ( .D(n12568), .CK(clk), .Q(img[964]), .QB(n31817) );
  DFFN img_reg_8__6__4_ ( .D(n12560), .CK(clk), .Q(img[972]), .QB(n31755) );
  DFFN img_reg_8__5__4_ ( .D(n12552), .CK(clk), .Q(img[980]), .QB(n31903) );
  DFFN img_reg_8__3__4_ ( .D(n12536), .CK(clk), .Q(img[996]), .QB(n31926) );
  DFFN img_reg_8__1__4_ ( .D(n12520), .CK(clk), .Q(img[1012]), .QB(n31950) );
  DFFN img_reg_6__6__2_ ( .D(n12302), .CK(clk), .Q(img[1226]), .QB(n30533) );
  DFFN img_reg_6__6__0_ ( .D(n12308), .CK(clk), .Q(img[1224]), .QB(n31641) );
  DFFN img_reg_5__6__2_ ( .D(n12178), .CK(clk), .Q(img[1354]), .QB(n30537) );
  DFFN img_reg_0__5__0_ ( .D(n11532), .CK(clk), .Q(img[2000]), .QB(n31633) );
  DFFN img_reg_6__0__0_ ( .D(n12260), .CK(clk), .Q(img[1272]), .QB(n31498) );
  DFFN img_reg_1__2__2_ ( .D(n11634), .CK(clk), .Q(img[1898]), .QB(n30558) );
  DFFN img_reg_1__0__2_ ( .D(n11618), .CK(clk), .Q(img[1914]), .QB(n30674) );
  DFFN img_reg_1__0__0_ ( .D(n11620), .CK(clk), .Q(img[1912]), .QB(n31506) );
  DFFN img_reg_6__1__2_ ( .D(n12266), .CK(clk), .Q(img[1266]), .QB(n30534) );
  DFFN img_reg_6__1__0_ ( .D(n12268), .CK(clk), .Q(img[1264]), .QB(n31642) );
  DFFN img_reg_5__1__2_ ( .D(n12134), .CK(clk), .Q(img[1394]), .QB(n30538) );
  DFFN img_reg_5__1__0_ ( .D(n12140), .CK(clk), .Q(img[1392]), .QB(n31646) );
  DFFN img_reg_2__3__2_ ( .D(n11770), .CK(clk), .Q(img[1762]), .QB(n30678) );
  DFFN img_reg_1__3__2_ ( .D(n11638), .CK(clk), .Q(img[1890]), .QB(n30670) );
  DFFN img_reg_1__3__0_ ( .D(n11644), .CK(clk), .Q(img[1888]), .QB(n31504) );
  DFFN img_reg_6__7__0_ ( .D(n12316), .CK(clk), .Q(img[1216]), .QB(n31500) );
  DFFN img_reg_3__7__0_ ( .D(n11932), .CK(clk), .Q(img[1600]), .QB(n31546) );
  DFFN img_reg_1__7__0_ ( .D(n11676), .CK(clk), .Q(img[1856]), .QB(n31508) );
  QDFFRBN img_size_reg_3_ ( .D(n13641), .CK(clk), .RB(n13805), .Q(img_size[3])
         );
  QDFFRBS rgb_value_reg_4_ ( .D(n11209), .CK(clk), .RB(n30035), .Q(
        rgb_value[4]) );
  DFFS img_reg_1__4__1_ ( .D(n11651), .CK(clk), .Q(img[1881]), .QB(n31039) );
  DFFS img_reg_5__10__7_ ( .D(n12205), .CK(clk), .Q(img[1327]), .QB(n30202) );
  DFFS img_reg_0__0__5_ ( .D(n11487), .CK(clk), .Q(img[2045]), .QB(n30827) );
  DFFS img_reg_4__2__2_ ( .D(n12014), .CK(clk), .Q(img[1514]), .QB(n30612) );
  DFFS img_reg_4__4__3_ ( .D(n12031), .CK(clk), .Q(img[1499]), .QB(n31459) );
  DFFS img_reg_0__0__3_ ( .D(n11489), .CK(clk), .Q(img[2043]), .QB(n31386) );
  DFFS img_reg_4__2__1_ ( .D(n12013), .CK(clk), .Q(img[1513]), .QB(n31140) );
  DFFS img_reg_4__0__7_ ( .D(n12003), .CK(clk), .Q(img[1535]), .QB(n30185) );
  DFFS img_reg_0__15__3_ ( .D(n11609), .CK(clk), .Q(img[1923]), .QB(n31385) );
  DFFS img_reg_5__15__2_ ( .D(n12246), .CK(clk), .Q(img[1282]), .QB(n30653) );
  DFFS img_reg_11__15__5_ ( .D(n13017), .CK(clk), .Q(img[517]), .QB(n30986) );
  DFFS img_reg_12__6__5_ ( .D(n13073), .CK(clk), .Q(img[461]), .QB(n30960) );
  DFFS img_reg_15__10__5_ ( .D(n13487), .CK(clk), .Q(img[45]), .QB(n30923) );
  DFFS img_reg_13__6__5_ ( .D(n13199), .CK(clk), .Q(img[333]), .QB(n30938) );
  DFFS img_reg_5__14__5_ ( .D(n12239), .CK(clk), .Q(img[1293]), .QB(n30951) );
  DFFS img_reg_4__10__3_ ( .D(n12079), .CK(clk), .Q(img[1451]), .QB(n31278) );
  DFFS img_reg_15__6__3_ ( .D(n13457), .CK(clk), .Q(img[75]), .QB(n31420) );
  DFFS img_reg_5__15__3_ ( .D(n12247), .CK(clk), .Q(img[1283]), .QB(n31340) );
  DFFS img_reg_13__12__3_ ( .D(n13249), .CK(clk), .Q(img[283]), .QB(n31489) );
  DFFS img_reg_1__14__3_ ( .D(n11729), .CK(clk), .Q(img[1803]), .QB(n31286) );
  DFFS img_reg_8__8__7_ ( .D(n12579), .CK(clk), .Q(img[959]), .QB(n30176) );
  DFFS img_reg_13__2__4_ ( .D(n13168), .CK(clk), .Q(img[364]), .QB(n31884) );
  DFFS img_reg_12__15__0_ ( .D(n13148), .CK(clk), .Q(img[384]), .QB(n31569) );
  DFFS img_reg_4__10__0_ ( .D(n12084), .CK(clk), .Q(img[1448]), .QB(n31593) );
  DFFS img_reg_15__14__2_ ( .D(n13522), .CK(clk), .Q(img[10]), .QB(n30531) );
  DFFS img_reg_7__15__0_ ( .D(n12508), .CK(clk), .Q(img[1024]), .QB(n31547) );
  DFFS img_reg_8__8__2_ ( .D(n12574), .CK(clk), .Q(img[954]), .QB(n30764) );
  DFFS img_reg_8__14__2_ ( .D(n12622), .CK(clk), .Q(img[906]), .QB(n30541) );
  DFFS img_reg_13__5__0_ ( .D(n13196), .CK(clk), .Q(img[336]), .QB(n31706) );
  DFFS img_reg_14__14__2_ ( .D(n13390), .CK(clk), .Q(img[138]), .QB(n30543) );
  DFFS img_reg_10__10__0_ ( .D(n12852), .CK(clk), .Q(img[680]), .QB(n31710) );
  DFFS img_reg_0__10__1_ ( .D(n11565), .CK(clk), .Q(img[1961]), .QB(n31180) );
  DFFS img_reg_9__9__1_ ( .D(n12709), .CK(clk), .Q(img[817]), .QB(n31225) );
  DFFS img_reg_7__11__1_ ( .D(n12469), .CK(clk), .Q(img[1057]), .QB(n31103) );
  DFFS img_reg_9__15__1_ ( .D(n12757), .CK(clk), .Q(img[769]), .QB(n31035) );
  DFFS img_reg_1__15__6_ ( .D(n11738), .CK(clk), .Q(img[1798]), .QB(n30312) );
  DFFS img_reg_2__8__1_ ( .D(n11805), .CK(clk), .Q(img[1721]), .QB(n31050) );
  DFFS img_reg_10__14__1_ ( .D(n12877), .CK(clk), .Q(img[649]), .QB(n31205) );
  DFFS img_reg_13__5__6_ ( .D(n13194), .CK(clk), .Q(img[342]), .QB(n30506) );
  DFFS img_reg_8__13__1_ ( .D(n12619), .CK(clk), .Q(img[913]), .QB(n31248) );
  DFFS img_reg_9__9__7_ ( .D(n12715), .CK(clk), .Q(img[823]), .QB(n30062) );
  DFFS img_reg_12__9__7_ ( .D(n13093), .CK(clk), .Q(img[439]), .QB(n30056) );
  DFFS img_reg_0__15__7_ ( .D(n11605), .CK(clk), .Q(img[1927]), .QB(n30158) );
  DFFS img_reg_13__10__7_ ( .D(n13229), .CK(clk), .Q(img[303]), .QB(n30232) );
  DFFS img_reg_11__15__4_ ( .D(n13016), .CK(clk), .Q(img[516]), .QB(n31974) );
  DFFS img_reg_12__9__4_ ( .D(n13096), .CK(clk), .Q(img[436]), .QB(n31760) );
  DFFS img_reg_5__15__4_ ( .D(n12248), .CK(clk), .Q(img[1284]), .QB(n31813) );
  DFFS img_reg_15__9__4_ ( .D(n13477), .CK(clk), .Q(img[52]), .QB(n31744) );
  DFFS img_reg_5__14__4_ ( .D(n12240), .CK(clk), .Q(img[1292]), .QB(n31750) );
  DFFS img_reg_10__8__4_ ( .D(n12832), .CK(clk), .Q(img[700]), .QB(n31830) );
  DFFS img_reg_10__6__5_ ( .D(n12817), .CK(clk), .Q(img[717]), .QB(n30943) );
  DFFS img_reg_10__4__6_ ( .D(n12802), .CK(clk), .Q(img[734]), .QB(n30467) );
  DFFS img_reg_10__2__7_ ( .D(n12787), .CK(clk), .Q(img[751]), .QB(n30219) );
  DFFS img_reg_10__1__0_ ( .D(n12780), .CK(clk), .Q(img[752]), .QB(n31661) );
  DFFS img_reg_0__11__1_ ( .D(n11579), .CK(clk), .Q(img[1953]), .QB(n31066) );
  DFFS img_reg_11__11__2_ ( .D(n12986), .CK(clk), .Q(img[546]), .QB(n30741) );
  DFFS img_reg_4__1__2_ ( .D(n12010), .CK(clk), .Q(img[1522]), .QB(n30550) );
  QDFFRBP i_col_reg_0_ ( .D(n13613), .CK(clk), .RB(n30034), .Q(i_col[0]) );
  QDFFRBS rgb_value_reg_15_ ( .D(n11220), .CK(clk), .RB(n30035), .Q(
        rgb_value[15]) );
  QDFFRBS rgb_value_reg_7_ ( .D(n11212), .CK(clk), .RB(n30035), .Q(
        rgb_value[7]) );
  QDFFRBS rgb_value_reg_6_ ( .D(n11211), .CK(clk), .RB(n30035), .Q(
        rgb_value[6]) );
  QDFFRBS rgb_value_reg_14_ ( .D(n11219), .CK(clk), .RB(n30035), .Q(
        rgb_value[14]) );
  QDFFRBS out_valid_reg ( .D(n31997), .CK(clk), .RB(n13805), .Q(out_valid) );
  QDFFRBS out_value_reg ( .D(N1330), .CK(clk), .RB(n13805), .Q(out_value) );
  QDFFRBS img_size_reg_4_ ( .D(n13640), .CK(clk), .RB(n13805), .Q(img_size[4])
         );
  QDFFS img_reg_9__8__0_ ( .D(n12708), .CK(clk), .Q(img[824]) );
  QDFFS img_reg_9__1__2_ ( .D(n12646), .CK(clk), .Q(img[882]) );
  QDFFS img_reg_9__1__3_ ( .D(n12647), .CK(clk), .Q(img[883]) );
  QDFFS img_reg_9__6__6_ ( .D(n12686), .CK(clk), .Q(img[846]) );
  QDFFS img_reg_9__2__7_ ( .D(n12653), .CK(clk), .Q(img[879]) );
  QDFFS img_reg_9__7__6_ ( .D(n12698), .CK(clk), .Q(img[838]) );
  QDFFS img_reg_9__4__6_ ( .D(n12670), .CK(clk), .Q(img[862]) );
  QDFFS img_reg_9__8__7_ ( .D(n12701), .CK(clk), .Q(img[831]) );
  QDFFS img_reg_9__0__6_ ( .D(n12638), .CK(clk), .Q(img[894]) );
  QDFFS img_reg_9__6__2_ ( .D(n12690), .CK(clk), .Q(img[842]) );
  QDFFS img_reg_9__3__1_ ( .D(n12661), .CK(clk), .Q(img[865]) );
  QDFFS img_reg_9__0__3_ ( .D(n12641), .CK(clk), .Q(img[891]) );
  QDFFS img_reg_9__5__6_ ( .D(n12682), .CK(clk), .Q(img[854]) );
  QDFFS img_reg_9__1__0_ ( .D(n12652), .CK(clk), .Q(img[880]) );
  QDFFS img_reg_9__2__6_ ( .D(n12654), .CK(clk), .Q(img[878]) );
  QDFFS img_reg_9__8__1_ ( .D(n12707), .CK(clk), .Q(img[825]) );
  QDFFS img_reg_9__8__6_ ( .D(n12702), .CK(clk), .Q(img[830]) );
  QDFFS img_reg_9__5__0_ ( .D(n12684), .CK(clk), .Q(img[848]) );
  QDFFS img_reg_9__7__0_ ( .D(n12700), .CK(clk), .Q(img[832]) );
  QDFFS img_reg_9__2__0_ ( .D(n12660), .CK(clk), .Q(img[872]) );
  QDFFS img_reg_9__5__2_ ( .D(n12678), .CK(clk), .Q(img[850]) );
  QDFFS img_reg_9__0__0_ ( .D(n12644), .CK(clk), .Q(img[888]) );
  QDFFS img_reg_9__8__2_ ( .D(n12706), .CK(clk), .Q(img[826]) );
  QDFFS img_reg_9__1__7_ ( .D(n12651), .CK(clk), .Q(img[887]) );
  QDFFS img_reg_9__1__6_ ( .D(n12650), .CK(clk), .Q(img[886]) );
  QDFFS img_reg_9__3__6_ ( .D(n12666), .CK(clk), .Q(img[870]) );
  QDFFS img_reg_9__4__0_ ( .D(n12676), .CK(clk), .Q(img[856]) );
  QDFFS img_reg_9__0__7_ ( .D(n12637), .CK(clk), .Q(img[895]) );
  QDFFS img_reg_9__6__7_ ( .D(n12685), .CK(clk), .Q(img[847]) );
  QDFFS img_reg_9__5__7_ ( .D(n12683), .CK(clk), .Q(img[855]) );
  QDFFS img_reg_9__3__0_ ( .D(n12668), .CK(clk), .Q(img[864]) );
  QDFFS img_reg_9__7__2_ ( .D(n12694), .CK(clk), .Q(img[834]) );
  QDFFS img_reg_9__8__3_ ( .D(n12705), .CK(clk), .Q(img[827]) );
  QDFFS img_reg_9__1__1_ ( .D(n12645), .CK(clk), .Q(img[881]) );
  QDFFS img_reg_9__3__7_ ( .D(n12667), .CK(clk), .Q(img[871]) );
  QDFFS img_reg_9__7__7_ ( .D(n12699), .CK(clk), .Q(img[839]) );
  QDFFS img_reg_9__4__2_ ( .D(n12674), .CK(clk), .Q(img[858]) );
  QDFFS img_reg_9__6__0_ ( .D(n12692), .CK(clk), .Q(img[840]) );
  QDFFS img_reg_9__2__1_ ( .D(n12659), .CK(clk), .Q(img[873]) );
  QDFFS img_reg_9__4__7_ ( .D(n12669), .CK(clk), .Q(img[863]) );
  QDFFS img_reg_9__2__2_ ( .D(n12658), .CK(clk), .Q(img[874]) );
  QDFFS img_reg_9__7__1_ ( .D(n12693), .CK(clk), .Q(img[833]) );
  QDFFS img_reg_9__4__1_ ( .D(n12675), .CK(clk), .Q(img[857]) );
  QDFFS img_reg_9__0__2_ ( .D(n12642), .CK(clk), .Q(img[890]) );
  QDFFS img_reg_9__5__1_ ( .D(n12677), .CK(clk), .Q(img[849]) );
  QDFFS img_reg_9__7__3_ ( .D(n12695), .CK(clk), .Q(img[835]) );
  QDFFS img_reg_12__0__7_ ( .D(n13027), .CK(clk), .Q(img[511]) );
  QDFFS img_reg_12__0__0_ ( .D(n13028), .CK(clk), .Q(img[504]) );
  QDFFS img_reg_12__0__6_ ( .D(n13026), .CK(clk), .Q(img[510]) );
  QDFFS img_reg_12__0__1_ ( .D(n13021), .CK(clk), .Q(img[505]) );
  QDFFS img_reg_12__0__2_ ( .D(n13022), .CK(clk), .Q(img[506]) );
  QDFFS img_reg_7__0__3_ ( .D(n12385), .CK(clk), .Q(img[1147]) );
  QDFFS img_reg_7__7__3_ ( .D(n12441), .CK(clk), .Q(img[1091]) );
  QDFFS img_reg_4__6__3_ ( .D(n12047), .CK(clk), .Q(img[1483]) );
  QDFFS img_reg_1__1__3_ ( .D(n11623), .CK(clk), .Q(img[1907]) );
  QDFFS img_reg_2__6__3_ ( .D(n11791), .CK(clk), .Q(img[1739]) );
  QDFFS img_reg_1__2__3_ ( .D(n11633), .CK(clk), .Q(img[1899]) );
  QDFFS img_reg_1__6__3_ ( .D(n11665), .CK(clk), .Q(img[1867]) );
  QDFFS img_reg_0__3__3_ ( .D(n11513), .CK(clk), .Q(img[2019]) );
  QDFFS img_reg_0__2__3_ ( .D(n11503), .CK(clk), .Q(img[2027]) );
  QDFFS img_reg_3__4__3_ ( .D(n11905), .CK(clk), .Q(img[1627]) );
  QDFFS img_reg_0__4__3_ ( .D(n11519), .CK(clk), .Q(img[2011]) );
  DFFS img_reg_4__5__7_ ( .D(n12037), .CK(clk), .Q(img[1495]), .QB(n30215) );
  DFFS img_reg_4__5__6_ ( .D(n12038), .CK(clk), .Q(img[1494]), .QB(n30488) );
  DFFS img_reg_4__5__1_ ( .D(n12043), .CK(clk), .Q(img[1489]), .QB(n31142) );
  DFFS img_reg_9__10__5_ ( .D(n12719), .CK(clk), .Q(img[813]), .QB(n30933) );
  DFFS img_reg_13__5__5_ ( .D(n13193), .CK(clk), .Q(img[341]), .QB(n30930) );
  DFFS img_reg_13__10__5_ ( .D(n13231), .CK(clk), .Q(img[301]), .QB(n30929) );
  DFFS img_reg_0__0__7_ ( .D(n13533), .CK(clk), .Q(img[2047]), .QB(n30159) );
  DFFS img_reg_1__4__6_ ( .D(n11646), .CK(clk), .Q(img[1886]), .QB(n30309) );
  DFFS img_reg_4__0__6_ ( .D(n12002), .CK(clk), .Q(img[1534]), .QB(n30303) );
  DFFS img_reg_3__4__1_ ( .D(n11907), .CK(clk), .Q(img[1625]), .QB(n31055) );
  DFFS img_reg_2__4__1_ ( .D(n11773), .CK(clk), .Q(img[1753]), .QB(n31047) );
  DFFS img_reg_0__4__7_ ( .D(n11523), .CK(clk), .Q(img[2015]), .QB(n30161) );
  DFFS img_reg_8__15__2_ ( .D(n12634), .CK(clk), .Q(img[898]), .QB(n30697) );
  DFFS img_reg_15__11__0_ ( .D(n13500), .CK(clk), .Q(img[32]), .QB(n31669) );
  DFFS img_reg_2__12__2_ ( .D(n11838), .CK(clk), .Q(img[1690]), .QB(n30677) );
  DFFS img_reg_7__8__2_ ( .D(n12450), .CK(clk), .Q(img[1082]), .QB(n30691) );
  DFFS img_reg_7__15__2_ ( .D(n12502), .CK(clk), .Q(img[1026]), .QB(n30693) );
  DFFS img_reg_3__8__2_ ( .D(n11938), .CK(clk), .Q(img[1594]), .QB(n30687) );
  DFFS img_reg_2__8__2_ ( .D(n11806), .CK(clk), .Q(img[1722]), .QB(n30679) );
  DFFS img_reg_3__12__2_ ( .D(n11970), .CK(clk), .Q(img[1562]), .QB(n30685) );
  DFFS img_reg_4__9__0_ ( .D(n12076), .CK(clk), .Q(img[1456]), .QB(n31656) );
  DFFS img_reg_3__15__2_ ( .D(n11990), .CK(clk), .Q(img[1538]), .QB(n30689) );
  DFFS img_reg_2__15__2_ ( .D(n11866), .CK(clk), .Q(img[1666]), .QB(n30681) );
  DFFS img_reg_13__1__0_ ( .D(n13164), .CK(clk), .Q(img[368]), .QB(n31652) );
  DFFS img_reg_0__4__4_ ( .D(n11520), .CK(clk), .Q(img[2012]), .QB(n31860) );
  DFFS img_reg_7__9__0_ ( .D(n12460), .CK(clk), .Q(img[1072]), .QB(n31663) );
  DFFS img_reg_3__11__2_ ( .D(n11958), .CK(clk), .Q(img[1570]), .QB(n30683) );
  DFFS img_reg_15__15__2_ ( .D(n13530), .CK(clk), .Q(img[2]), .QB(n30695) );
  DFFS img_reg_4__9__3_ ( .D(n12073), .CK(clk), .Q(img[1459]), .QB(n31409) );
  DFFS img_reg_15__9__3_ ( .D(n13481), .CK(clk), .Q(img[51]), .QB(n31419) );
  DFFS img_reg_13__1__3_ ( .D(n13159), .CK(clk), .Q(img[371]), .QB(n31405) );
  DFFS img_reg_15__1__1_ ( .D(n13413), .CK(clk), .Q(img[113]), .QB(n31190) );
  DFFS img_reg_15__4__6_ ( .D(n13438), .CK(clk), .Q(img[94]), .QB(n30456) );
  DFFS img_reg_7__12__6_ ( .D(n12478), .CK(clk), .Q(img[1054]), .QB(n30437) );
  DFFS img_reg_15__9__6_ ( .D(n13479), .CK(clk), .Q(img[54]), .QB(n30440) );
  DFFS img_reg_13__6__6_ ( .D(n13198), .CK(clk), .Q(img[334]), .QB(n30447) );
  DFFS img_reg_13__9__6_ ( .D(n13226), .CK(clk), .Q(img[310]), .QB(n30446) );
  DFFS img_reg_6__10__7_ ( .D(n12339), .CK(clk), .Q(img[1199]), .QB(n30198) );
  DFFS img_reg_4__13__7_ ( .D(n12101), .CK(clk), .Q(img[1431]), .QB(n30217) );
  DFFS img_reg_6__13__7_ ( .D(n12357), .CK(clk), .Q(img[1175]), .QB(n30201) );
  DFFS img_reg_13__13__7_ ( .D(n13259), .CK(clk), .Q(img[279]), .QB(n30211) );
  DFFS img_reg_15__13__7_ ( .D(n13515), .CK(clk), .Q(img[23]), .QB(n30197) );
  DFFS img_reg_13__2__7_ ( .D(n13165), .CK(clk), .Q(img[367]), .QB(n30210) );
  DFFS img_reg_11__13__7_ ( .D(n13003), .CK(clk), .Q(img[535]), .QB(n30195) );
  DFFS img_reg_7__13__1_ ( .D(n12491), .CK(clk), .Q(img[1041]), .QB(n31170) );
  DFFS img_reg_9__9__6_ ( .D(n12714), .CK(clk), .Q(img[822]), .QB(n30450) );
  DFFS img_reg_3__9__1_ ( .D(n11941), .CK(clk), .Q(img[1585]), .QB(n31162) );
  DFFS img_reg_15__14__1_ ( .D(n13523), .CK(clk), .Q(img[9]), .QB(n31189) );
  DFFS img_reg_2__4__5_ ( .D(n11777), .CK(clk), .Q(img[1757]), .QB(n30811) );
  DFFS img_reg_9__10__4_ ( .D(n12720), .CK(clk), .Q(img[812]), .QB(n31910) );
  DFFS img_reg_4__1__5_ ( .D(n12007), .CK(clk), .Q(img[1525]), .QB(n30962) );
  DFFS img_reg_4__0__5_ ( .D(n12001), .CK(clk), .Q(img[1533]), .QB(n30909) );
  DFFS img_reg_0__4__5_ ( .D(n11521), .CK(clk), .Q(img[2013]), .QB(n30829) );
  DFFS img_reg_3__4__5_ ( .D(n11903), .CK(clk), .Q(img[1629]), .QB(n30818) );
  DFFS img_reg_7__11__4_ ( .D(n12472), .CK(clk), .Q(img[1060]), .QB(n31915) );
  DFFS img_reg_4__4__5_ ( .D(n12033), .CK(clk), .Q(img[1501]), .QB(n30795) );
  DFFS img_reg_4__2__5_ ( .D(n12017), .CK(clk), .Q(img[1517]), .QB(n30854) );
  DFFS img_reg_13__5__4_ ( .D(n13192), .CK(clk), .Q(img[340]), .QB(n31907) );
  DFFS img_reg_13__3__4_ ( .D(n13176), .CK(clk), .Q(img[356]), .QB(n31914) );
  DFFS img_reg_13__10__4_ ( .D(n13232), .CK(clk), .Q(img[300]), .QB(n31906) );
  DFFS img_reg_3__4__0_ ( .D(n11908), .CK(clk), .Q(img[1624]), .QB(n31540) );
  DFFS img_reg_2__4__0_ ( .D(n11780), .CK(clk), .Q(img[1752]), .QB(n31532) );
  DFFS img_reg_4__4__0_ ( .D(n12036), .CK(clk), .Q(img[1496]), .QB(n31690) );
  DFFS img_reg_4__2__0_ ( .D(n12020), .CK(clk), .Q(img[1512]), .QB(n31596) );
  DFFS img_reg_4__0__2_ ( .D(n11998), .CK(clk), .Q(img[1530]), .QB(n30663) );
  DFFS img_reg_4__0__0_ ( .D(n12004), .CK(clk), .Q(img[1528]), .QB(n31512) );
  DFFS img_reg_0__4__0_ ( .D(n11524), .CK(clk), .Q(img[2008]), .QB(n31552) );
  DFFS img_reg_3__4__2_ ( .D(n11906), .CK(clk), .Q(img[1626]), .QB(n30684) );
  DFFS img_reg_0__4__2_ ( .D(n11518), .CK(clk), .Q(img[2010]), .QB(n30642) );
  DFFS img_reg_4__4__2_ ( .D(n12030), .CK(clk), .Q(img[1498]), .QB(n30733) );
  DFFS img_reg_4__3__2_ ( .D(n12026), .CK(clk), .Q(img[1506]), .QB(n30731) );
  DFFS img_reg_4__3__0_ ( .D(n12028), .CK(clk), .Q(img[1504]), .QB(n31688) );
  DFFS img_reg_4__1__0_ ( .D(n12012), .CK(clk), .Q(img[1520]), .QB(n31658) );
  DFFS img_reg_0__0__2_ ( .D(n11490), .CK(clk), .Q(img[2042]), .QB(n30648) );
  DFFS img_reg_0__0__0_ ( .D(n11492), .CK(clk), .Q(img[2040]), .QB(n31556) );
  DFFS img_reg_2__4__3_ ( .D(n11775), .CK(clk), .Q(img[1755]), .QB(n31367) );
  DFFS img_reg_1__4__3_ ( .D(n11649), .CK(clk), .Q(img[1883]), .QB(n31359) );
  DFFS img_reg_4__3__3_ ( .D(n12025), .CK(clk), .Q(img[1507]), .QB(n31457) );
  DFFS img_reg_4__2__3_ ( .D(n12015), .CK(clk), .Q(img[1515]), .QB(n31279) );
  DFFS img_reg_4__1__3_ ( .D(n12009), .CK(clk), .Q(img[1523]), .QB(n31410) );
  DFFS img_reg_4__0__3_ ( .D(n11999), .CK(clk), .Q(img[1531]), .QB(n31353) );
  DFFS img_reg_3__4__6_ ( .D(n11902), .CK(clk), .Q(img[1630]), .QB(n30325) );
  DFFS img_reg_2__4__6_ ( .D(n11778), .CK(clk), .Q(img[1758]), .QB(n30317) );
  DFFS img_reg_4__4__6_ ( .D(n12034), .CK(clk), .Q(img[1502]), .QB(n30428) );
  DFFS img_reg_4__4__1_ ( .D(n12029), .CK(clk), .Q(img[1497]), .QB(n31095) );
  DFFS img_reg_4__0__1_ ( .D(n11997), .CK(clk), .Q(img[1529]), .QB(n31032) );
  DFFS img_reg_0__4__6_ ( .D(n11522), .CK(clk), .Q(img[2014]), .QB(n30337) );
  DFFS img_reg_0__4__1_ ( .D(n11517), .CK(clk), .Q(img[2009]), .QB(n31067) );
  DFFS img_reg_4__3__6_ ( .D(n12022), .CK(clk), .Q(img[1510]), .QB(n30429) );
  DFFS img_reg_4__3__1_ ( .D(n12027), .CK(clk), .Q(img[1505]), .QB(n31094) );
  DFFS img_reg_4__1__6_ ( .D(n12006), .CK(clk), .Q(img[1526]), .QB(n30367) );
  DFFS img_reg_4__2__6_ ( .D(n12018), .CK(clk), .Q(img[1518]), .QB(n30487) );
  DFFS img_reg_4__1__1_ ( .D(n12011), .CK(clk), .Q(img[1521]), .QB(n31204) );
  DFFS img_reg_3__4__7_ ( .D(n11901), .CK(clk), .Q(img[1631]), .QB(n30149) );
  DFFS img_reg_2__4__7_ ( .D(n11779), .CK(clk), .Q(img[1759]), .QB(n30141) );
  DFFS img_reg_1__4__7_ ( .D(n11645), .CK(clk), .Q(img[1887]), .QB(n30133) );
  DFFS img_reg_4__4__7_ ( .D(n12035), .CK(clk), .Q(img[1503]), .QB(n30122) );
  DFFS img_reg_4__3__7_ ( .D(n12021), .CK(clk), .Q(img[1511]), .QB(n30123) );
  DFFS img_reg_4__1__7_ ( .D(n12005), .CK(clk), .Q(img[1527]), .QB(n30059) );
  DFFS img_reg_4__2__7_ ( .D(n12019), .CK(clk), .Q(img[1519]), .QB(n30216) );
  DFFS img_reg_10__14__3_ ( .D(n12879), .CK(clk), .Q(img[651]), .QB(n31414) );
  DFFS img_reg_9__14__1_ ( .D(n12755), .CK(clk), .Q(img[777]), .QB(n31186) );
  DFFS img_reg_9__14__0_ ( .D(n12756), .CK(clk), .Q(img[776]), .QB(n31660) );
  DFFS img_reg_8__14__3_ ( .D(n12623), .CK(clk), .Q(img[907]), .QB(n31402) );
  DFFS img_reg_8__14__0_ ( .D(n12628), .CK(clk), .Q(img[904]), .QB(n31649) );
  DFFS img_reg_0__0__1_ ( .D(n11491), .CK(clk), .Q(img[2041]), .QB(n31072) );
  DFFS img_reg_0__0__6_ ( .D(n11486), .CK(clk), .Q(img[2046]), .QB(n30341) );
  DFFS img_reg_3__4__4_ ( .D(n11904), .CK(clk), .Q(img[1628]), .QB(n31848) );
  DFFS img_reg_2__4__4_ ( .D(n11776), .CK(clk), .Q(img[1756]), .QB(n31840) );
  DFFS img_reg_1__4__4_ ( .D(n11648), .CK(clk), .Q(img[1884]), .QB(n31832) );
  DFFS img_reg_4__4__4_ ( .D(n12032), .CK(clk), .Q(img[1500]), .QB(n31934) );
  DFFS img_reg_4__3__4_ ( .D(n12024), .CK(clk), .Q(img[1508]), .QB(n31936) );
  DFFS img_reg_4__1__4_ ( .D(n12008), .CK(clk), .Q(img[1524]), .QB(n31763) );
  DFFS img_reg_4__0__4_ ( .D(n12000), .CK(clk), .Q(img[1532]), .QB(n31826) );
  DFFS img_reg_4__2__4_ ( .D(n12016), .CK(clk), .Q(img[1516]), .QB(n31890) );
  DFFS img_reg_0__0__4_ ( .D(n11488), .CK(clk), .Q(img[2044]), .QB(n31864) );
  DFFS img_reg_9__8__5_ ( .D(n12703), .CK(clk), .Q(img[829]), .QB(n30912) );
  DFFS img_reg_7__15__5_ ( .D(n12505), .CK(clk), .Q(img[1029]), .QB(n30913) );
  DFFS img_reg_6__15__5_ ( .D(n12375), .CK(clk), .Q(img[1157]), .QB(n30898) );
  DFFS img_reg_5__15__5_ ( .D(n12249), .CK(clk), .Q(img[1285]), .QB(n30900) );
  DFFS img_reg_4__15__5_ ( .D(n12119), .CK(clk), .Q(img[1413]), .QB(n30908) );
  DFFS img_reg_8__8__5_ ( .D(n12577), .CK(clk), .Q(img[957]), .QB(n30902) );
  DFFS img_reg_4__8__5_ ( .D(n12065), .CK(clk), .Q(img[1469]), .QB(n30910) );
  DFFS img_reg_7__8__5_ ( .D(n12447), .CK(clk), .Q(img[1085]), .QB(n30915) );
  DFFS img_reg_5__8__5_ ( .D(n12191), .CK(clk), .Q(img[1341]), .QB(n30901) );
  DFFS img_reg_13__8__5_ ( .D(n13215), .CK(clk), .Q(img[317]), .QB(n30904) );
  DFFS img_reg_13__7__5_ ( .D(n13209), .CK(clk), .Q(img[325]), .QB(n30905) );
  DFFS img_reg_3__11__3_ ( .D(n11959), .CK(clk), .Q(img[1571]), .QB(n31374) );
  DFFS img_reg_8__6__6_ ( .D(n12562), .CK(clk), .Q(img[974]), .QB(n30443) );
  DFFS img_reg_8__2__7_ ( .D(n12531), .CK(clk), .Q(img[1007]), .QB(n30206) );
  DFFS img_reg_8__1__3_ ( .D(n12521), .CK(clk), .Q(img[1011]), .QB(n31401) );
  DFFS img_reg_15__14__3_ ( .D(n13521), .CK(clk), .Q(img[11]), .QB(n31392) );
  DFFS img_reg_7__15__3_ ( .D(n12503), .CK(clk), .Q(img[1027]), .QB(n31381) );
  DFFS img_reg_3__15__3_ ( .D(n11991), .CK(clk), .Q(img[1539]), .QB(n31377) );
  DFFS img_reg_2__15__3_ ( .D(n11865), .CK(clk), .Q(img[1667]), .QB(n31370) );
  DFFS img_reg_6__9__3_ ( .D(n12329), .CK(clk), .Q(img[1203]), .QB(n31393) );
  DFFS img_reg_7__8__3_ ( .D(n12449), .CK(clk), .Q(img[1083]), .QB(n31382) );
  DFFS img_reg_3__8__3_ ( .D(n11937), .CK(clk), .Q(img[1595]), .QB(n31379) );
  DFFS img_reg_2__8__3_ ( .D(n11807), .CK(clk), .Q(img[1723]), .QB(n31372) );
  DFFS img_reg_11__14__3_ ( .D(n13009), .CK(clk), .Q(img[523]), .QB(n31390) );
  DFFS img_reg_6__14__3_ ( .D(n12367), .CK(clk), .Q(img[1163]), .QB(n31396) );
  DFFS img_reg_1__11__2_ ( .D(n11702), .CK(clk), .Q(img[1826]), .QB(n30667) );
  DFFS img_reg_12__15__2_ ( .D(n13146), .CK(clk), .Q(img[386]), .QB(n30659) );
  DFFS img_reg_11__15__2_ ( .D(n13014), .CK(clk), .Q(img[514]), .QB(n30649) );
  DFFS img_reg_3__9__0_ ( .D(n11948), .CK(clk), .Q(img[1584]), .QB(n31616) );
  DFFS img_reg_15__14__0_ ( .D(n13524), .CK(clk), .Q(img[8]), .QB(n31639) );
  DFFS img_reg_1__12__2_ ( .D(n11714), .CK(clk), .Q(img[1818]), .QB(n30669) );
  DFFS img_reg_13__15__2_ ( .D(n13270), .CK(clk), .Q(img[258]), .QB(n30657) );
  DFFS img_reg_10__15__2_ ( .D(n12890), .CK(clk), .Q(img[642]), .QB(n30665) );
  DFFS img_reg_9__15__2_ ( .D(n12758), .CK(clk), .Q(img[770]), .QB(n30664) );
  DFFS img_reg_4__15__2_ ( .D(n12122), .CK(clk), .Q(img[1410]), .QB(n30662) );
  DFFS img_reg_1__15__2_ ( .D(n11734), .CK(clk), .Q(img[1794]), .QB(n30673) );
  DFFS img_reg_0__15__2_ ( .D(n11610), .CK(clk), .Q(img[1922]), .QB(n30647) );
  DFFS img_reg_6__9__0_ ( .D(n12332), .CK(clk), .Q(img[1200]), .QB(n31640) );
  DFFS img_reg_4__8__2_ ( .D(n12062), .CK(clk), .Q(img[1466]), .QB(n30660) );
  DFFS img_reg_5__8__2_ ( .D(n12194), .CK(clk), .Q(img[1338]), .QB(n30651) );
  DFFS img_reg_11__14__0_ ( .D(n13012), .CK(clk), .Q(img[520]), .QB(n31637) );
  DFFS img_reg_6__14__0_ ( .D(n12372), .CK(clk), .Q(img[1160]), .QB(n31643) );
  DFFS img_reg_4__10__7_ ( .D(n12083), .CK(clk), .Q(img[1455]), .QB(n30214) );
  DFFS img_reg_13__0__2_ ( .D(n13154), .CK(clk), .Q(img[378]), .QB(n30658) );
  DFFS img_reg_8__13__7_ ( .D(n12613), .CK(clk), .Q(img[919]), .QB(n30207) );
  DFFS img_reg_1__11__5_ ( .D(n11705), .CK(clk), .Q(img[1829]), .QB(n30803) );
  DFFS img_reg_12__15__5_ ( .D(n13143), .CK(clk), .Q(img[389]), .QB(n30992) );
  DFFS img_reg_3__9__5_ ( .D(n11945), .CK(clk), .Q(img[1589]), .QB(n30875) );
  DFFS img_reg_9__9__5_ ( .D(n12713), .CK(clk), .Q(img[821]), .QB(n30965) );
  DFFS img_reg_5__10__5_ ( .D(n12207), .CK(clk), .Q(img[1325]), .QB(n30840) );
  DFFS img_reg_9__6__5_ ( .D(n12687), .CK(clk), .Q(img[845]), .QB(n30966) );
  DFFS img_reg_9__5__5_ ( .D(n12681), .CK(clk), .Q(img[853]), .QB(n30934) );
  DFFS img_reg_9__4__5_ ( .D(n12671), .CK(clk), .Q(img[861]), .QB(n31008) );
  DFFS img_reg_4__10__5_ ( .D(n12081), .CK(clk), .Q(img[1453]), .QB(n30852) );
  DFFS img_reg_15__15__5_ ( .D(n13527), .CK(clk), .Q(img[5]), .QB(n30988) );
  DFFS img_reg_7__11__5_ ( .D(n12473), .CK(clk), .Q(img[1061]), .QB(n30820) );
  DFFS img_reg_3__11__5_ ( .D(n11961), .CK(clk), .Q(img[1573]), .QB(n30817) );
  DFFS img_reg_10__11__5_ ( .D(n12855), .CK(clk), .Q(img[677]), .QB(n31009) );
  DFFS img_reg_9__11__5_ ( .D(n12729), .CK(clk), .Q(img[805]), .QB(n31007) );
  DFFS img_reg_4__11__5_ ( .D(n12087), .CK(clk), .Q(img[1445]), .QB(n30794) );
  DFFS img_reg_12__9__5_ ( .D(n13095), .CK(clk), .Q(img[437]), .QB(n30959) );
  DFFS img_reg_15__14__5_ ( .D(n13519), .CK(clk), .Q(img[13]), .QB(n30969) );
  DFFS img_reg_15__6__5_ ( .D(n13455), .CK(clk), .Q(img[77]), .QB(n30947) );
  DFFS img_reg_7__12__5_ ( .D(n12479), .CK(clk), .Q(img[1053]), .QB(n30822) );
  DFFS img_reg_6__10__5_ ( .D(n12337), .CK(clk), .Q(img[1197]), .QB(n30836) );
  DFFS img_reg_8__6__5_ ( .D(n12561), .CK(clk), .Q(img[973]), .QB(n30956) );
  DFFS img_reg_8__0__5_ ( .D(n12513), .CK(clk), .Q(img[1021]), .QB(n30991) );
  DFFS img_reg_6__13__5_ ( .D(n12359), .CK(clk), .Q(img[1173]), .QB(n30839) );
  DFFS img_reg_4__13__5_ ( .D(n12103), .CK(clk), .Q(img[1429]), .QB(n30855) );
  DFFS img_reg_13__15__5_ ( .D(n13273), .CK(clk), .Q(img[261]), .QB(n30984) );
  DFFS img_reg_10__15__5_ ( .D(n12887), .CK(clk), .Q(img[645]), .QB(n30994) );
  DFFS img_reg_9__15__5_ ( .D(n12761), .CK(clk), .Q(img[773]), .QB(n30993) );
  DFFS img_reg_8__15__5_ ( .D(n12631), .CK(clk), .Q(img[901]), .QB(n30990) );
  DFFS img_reg_3__15__5_ ( .D(n11993), .CK(clk), .Q(img[1541]), .QB(n30815) );
  DFFS img_reg_2__15__5_ ( .D(n11863), .CK(clk), .Q(img[1669]), .QB(n30808) );
  DFFS img_reg_1__15__5_ ( .D(n11737), .CK(clk), .Q(img[1797]), .QB(n30801) );
  DFFS img_reg_0__15__5_ ( .D(n11607), .CK(clk), .Q(img[1925]), .QB(n30826) );
  DFFS img_reg_6__9__5_ ( .D(n12327), .CK(clk), .Q(img[1205]), .QB(n30950) );
  DFFS img_reg_4__9__5_ ( .D(n12071), .CK(clk), .Q(img[1461]), .QB(n30963) );
  DFFS img_reg_13__13__5_ ( .D(n13257), .CK(clk), .Q(img[277]), .QB(n30849) );
  DFFS img_reg_15__13__5_ ( .D(n13513), .CK(clk), .Q(img[21]), .QB(n30835) );
  DFFS img_reg_3__8__5_ ( .D(n11935), .CK(clk), .Q(img[1597]), .QB(n30814) );
  DFFS img_reg_2__8__5_ ( .D(n11809), .CK(clk), .Q(img[1725]), .QB(n30806) );
  DFFS img_reg_15__9__5_ ( .D(n13478), .CK(clk), .Q(img[53]), .QB(n30946) );
  DFFS img_reg_11__14__5_ ( .D(n13007), .CK(clk), .Q(img[525]), .QB(n30971) );
  DFFS img_reg_10__14__5_ ( .D(n12881), .CK(clk), .Q(img[653]), .QB(n30980) );
  DFFS img_reg_9__14__5_ ( .D(n12751), .CK(clk), .Q(img[781]), .QB(n30979) );
  DFFS img_reg_8__14__5_ ( .D(n12625), .CK(clk), .Q(img[909]), .QB(n30973) );
  DFFS img_reg_6__14__5_ ( .D(n12369), .CK(clk), .Q(img[1165]), .QB(n30948) );
  DFFS img_reg_13__12__5_ ( .D(n13247), .CK(clk), .Q(img[285]), .QB(n30790) );
  DFFS img_reg_13__11__5_ ( .D(n13241), .CK(clk), .Q(img[293]), .QB(n31003) );
  DFFS img_reg_13__4__5_ ( .D(n13183), .CK(clk), .Q(img[349]), .QB(n31004) );
  DFFS img_reg_13__3__5_ ( .D(n13177), .CK(clk), .Q(img[357]), .QB(n30791) );
  DFFS img_reg_13__2__5_ ( .D(n13167), .CK(clk), .Q(img[365]), .QB(n30848) );
  DFFS img_reg_13__1__5_ ( .D(n13161), .CK(clk), .Q(img[373]), .QB(n30978) );
  DFFS img_reg_13__0__5_ ( .D(n13151), .CK(clk), .Q(img[381]), .QB(n30985) );
  DFFS img_reg_10__13__5_ ( .D(n12871), .CK(clk), .Q(img[661]), .QB(n30858) );
  DFFS img_reg_9__13__5_ ( .D(n12745), .CK(clk), .Q(img[789]), .QB(n30856) );
  DFFS img_reg_8__13__5_ ( .D(n12615), .CK(clk), .Q(img[917]), .QB(n30845) );
  DFFS img_reg_12__13__5_ ( .D(n13127), .CK(clk), .Q(img[405]), .QB(n30851) );
  DFFS img_reg_11__13__5_ ( .D(n13001), .CK(clk), .Q(img[533]), .QB(n30833) );
  DFFS img_reg_13__9__5_ ( .D(n13225), .CK(clk), .Q(img[309]), .QB(n30937) );
  DFFS img_reg_14__14__5_ ( .D(n13393), .CK(clk), .Q(img[141]), .QB(n30975) );
  DFFS img_reg_14__14__3_ ( .D(n13391), .CK(clk), .Q(img[139]), .QB(n31404) );
  DFFS img_reg_14__14__0_ ( .D(n13396), .CK(clk), .Q(img[136]), .QB(n31651) );
  DFFS img_reg_5__14__3_ ( .D(n12241), .CK(clk), .Q(img[1291]), .QB(n31400) );
  DFFS img_reg_5__14__0_ ( .D(n12244), .CK(clk), .Q(img[1288]), .QB(n31647) );
  DFFS img_reg_3__14__5_ ( .D(n11983), .CK(clk), .Q(img[1549]), .QB(n30877) );
  DFFS img_reg_3__14__1_ ( .D(n11987), .CK(clk), .Q(img[1545]), .QB(n31164) );
  DFFS img_reg_3__14__0_ ( .D(n11988), .CK(clk), .Q(img[1544]), .QB(n31618) );
  DFFS img_reg_1__14__5_ ( .D(n11727), .CK(clk), .Q(img[1805]), .QB(n30861) );
  DFFS img_reg_12__14__3_ ( .D(n13135), .CK(clk), .Q(img[395]), .QB(n31408) );
  DFFS img_reg_12__14__0_ ( .D(n13140), .CK(clk), .Q(img[392]), .QB(n31655) );
  DFFS img_reg_8__9__6_ ( .D(n12582), .CK(clk), .Q(img[950]), .QB(n30442) );
  DFFS img_reg_8__9__5_ ( .D(n12583), .CK(clk), .Q(img[949]), .QB(n30955) );
  DFFS img_reg_1__9__1_ ( .D(n11685), .CK(clk), .Q(img[1841]), .QB(n31146) );
  DFFS img_reg_5__10__1_ ( .D(n12211), .CK(clk), .Q(img[1321]), .QB(n31129) );
  DFFS img_reg_9__10__1_ ( .D(n12723), .CK(clk), .Q(img[809]), .QB(n31143) );
  DFFS img_reg_4__10__1_ ( .D(n12077), .CK(clk), .Q(img[1449]), .QB(n31141) );
  DFFS img_reg_7__13__3_ ( .D(n12486), .CK(clk), .Q(img[1043]), .QB(n31308) );
  DFFS img_reg_2__13__3_ ( .D(n11849), .CK(clk), .Q(img[1683]), .QB(n31296) );
  DFFS img_reg_1__13__3_ ( .D(n11719), .CK(clk), .Q(img[1811]), .QB(n31289) );
  DFFS img_reg_1__11__3_ ( .D(n11703), .CK(clk), .Q(img[1827]), .QB(n31358) );
  DFFS img_reg_4__11__6_ ( .D(n12086), .CK(clk), .Q(img[1446]), .QB(n30427) );
  DFFS img_reg_12__15__3_ ( .D(n13145), .CK(clk), .Q(img[387]), .QB(n31466) );
  DFFS img_reg_11__15__3_ ( .D(n13015), .CK(clk), .Q(img[515]), .QB(n31468) );
  DFFS img_reg_3__9__3_ ( .D(n11943), .CK(clk), .Q(img[1587]), .QB(n31297) );
  DFFS img_reg_9__9__3_ ( .D(n12711), .CK(clk), .Q(img[819]), .QB(n31427) );
  DFFS img_reg_8__9__3_ ( .D(n12585), .CK(clk), .Q(img[947]), .QB(n31421) );
  DFFS img_reg_5__10__3_ ( .D(n12209), .CK(clk), .Q(img[1323]), .QB(n31266) );
  DFFS img_reg_9__6__3_ ( .D(n12689), .CK(clk), .Q(img[843]), .QB(n31428) );
  DFFS img_reg_9__5__3_ ( .D(n12679), .CK(clk), .Q(img[851]), .QB(n31328) );
  DFFS img_reg_9__4__3_ ( .D(n12673), .CK(clk), .Q(img[859]), .QB(n31465) );
  DFFS img_reg_9__3__3_ ( .D(n12663), .CK(clk), .Q(img[867]), .QB(n31494) );
  DFFS img_reg_9__2__3_ ( .D(n12657), .CK(clk), .Q(img[875]), .QB(n31281) );
  DFFS img_reg_9__10__3_ ( .D(n12721), .CK(clk), .Q(img[811]), .QB(n31329) );
  DFFS img_reg_15__15__3_ ( .D(n13529), .CK(clk), .Q(img[3]), .QB(n31470) );
  DFFS img_reg_7__11__3_ ( .D(n12471), .CK(clk), .Q(img[1059]), .QB(n31439) );
  DFFS img_reg_2__14__1_ ( .D(n11853), .CK(clk), .Q(img[1673]), .QB(n31156) );
  DFFS img_reg_12__10__1_ ( .D(n13101), .CK(clk), .Q(img[425]), .QB(n31137) );
  DFFS img_reg_15__12__6_ ( .D(n13502), .CK(clk), .Q(img[30]), .QB(n30410) );
  DFFS img_reg_12__12__6_ ( .D(n13122), .CK(clk), .Q(img[414]), .QB(n30426) );
  DFFS img_reg_15__3__6_ ( .D(n13434), .CK(clk), .Q(img[102]), .QB(n30409) );
  DFFS img_reg_11__12__6_ ( .D(n12990), .CK(clk), .Q(img[542]), .QB(n30408) );
  DFFS img_reg_10__12__6_ ( .D(n12866), .CK(clk), .Q(img[670]), .QB(n30433) );
  DFFS img_reg_9__12__6_ ( .D(n12734), .CK(clk), .Q(img[798]), .QB(n30431) );
  DFFS img_reg_8__12__6_ ( .D(n12610), .CK(clk), .Q(img[926]), .QB(n30420) );
  DFFS img_reg_6__12__6_ ( .D(n12354), .CK(clk), .Q(img[1182]), .QB(n30414) );
  DFFS img_reg_10__11__3_ ( .D(n12857), .CK(clk), .Q(img[675]), .QB(n31460) );
  DFFS img_reg_9__11__3_ ( .D(n12727), .CK(clk), .Q(img[803]), .QB(n31464) );
  DFFS img_reg_4__11__3_ ( .D(n12089), .CK(clk), .Q(img[1443]), .QB(n31458) );
  DFFS img_reg_8__5__1_ ( .D(n12555), .CK(clk), .Q(img[977]), .QB(n31132) );
  DFFS img_reg_8__3__6_ ( .D(n12534), .CK(clk), .Q(img[998]), .QB(n30419) );
  DFFS img_reg_12__9__3_ ( .D(n13097), .CK(clk), .Q(img[435]), .QB(n31431) );
  DFFS img_reg_12__6__3_ ( .D(n13071), .CK(clk), .Q(img[459]), .QB(n31432) );
  DFFS img_reg_4__13__1_ ( .D(n12107), .CK(clk), .Q(img[1425]), .QB(n31139) );
  DFFS img_reg_7__14__3_ ( .D(n12497), .CK(clk), .Q(img[1035]), .QB(n31418) );
  DFFS img_reg_2__14__3_ ( .D(n11855), .CK(clk), .Q(img[1675]), .QB(n31291) );
  DFFS img_reg_12__10__3_ ( .D(n13103), .CK(clk), .Q(img[427]), .QB(n31327) );
  DFFS img_reg_15__12__3_ ( .D(n13505), .CK(clk), .Q(img[27]), .QB(n31483) );
  DFFS img_reg_15__11__3_ ( .D(n13495), .CK(clk), .Q(img[35]), .QB(n31442) );
  DFFS img_reg_12__12__3_ ( .D(n13119), .CK(clk), .Q(img[411]), .QB(n31491) );
  DFFS img_reg_7__12__3_ ( .D(n12481), .CK(clk), .Q(img[1051]), .QB(n31437) );
  DFFS img_reg_15__4__3_ ( .D(n13441), .CK(clk), .Q(img[91]), .QB(n31443) );
  DFFS img_reg_15__3__3_ ( .D(n13431), .CK(clk), .Q(img[99]), .QB(n31484) );
  DFFS img_reg_11__12__3_ ( .D(n12993), .CK(clk), .Q(img[539]), .QB(n31481) );
  DFFS img_reg_10__12__3_ ( .D(n12863), .CK(clk), .Q(img[667]), .QB(n31495) );
  DFFS img_reg_9__12__3_ ( .D(n12737), .CK(clk), .Q(img[795]), .QB(n31493) );
  DFFS img_reg_8__12__3_ ( .D(n12607), .CK(clk), .Q(img[923]), .QB(n31485) );
  DFFS img_reg_6__10__3_ ( .D(n12335), .CK(clk), .Q(img[1195]), .QB(n31262) );
  DFFS img_reg_8__6__3_ ( .D(n12559), .CK(clk), .Q(img[971]), .QB(n31422) );
  DFFS img_reg_8__5__3_ ( .D(n12553), .CK(clk), .Q(img[979]), .QB(n31320) );
  DFFS img_reg_8__3__3_ ( .D(n12537), .CK(clk), .Q(img[995]), .QB(n31486) );
  DFFS img_reg_8__2__3_ ( .D(n12527), .CK(clk), .Q(img[1003]), .QB(n31270) );
  DFFS img_reg_6__13__3_ ( .D(n12361), .CK(clk), .Q(img[1171]), .QB(n31265) );
  DFFS img_reg_4__13__3_ ( .D(n12105), .CK(clk), .Q(img[1427]), .QB(n31280) );
  DFFS img_reg_13__15__3_ ( .D(n13271), .CK(clk), .Q(img[259]), .QB(n31476) );
  DFFS img_reg_10__15__3_ ( .D(n12889), .CK(clk), .Q(img[643]), .QB(n31479) );
  DFFS img_reg_9__15__3_ ( .D(n12759), .CK(clk), .Q(img[771]), .QB(n31478) );
  DFFS img_reg_8__15__3_ ( .D(n12633), .CK(clk), .Q(img[899]), .QB(n31472) );
  DFFS img_reg_6__15__3_ ( .D(n12377), .CK(clk), .Q(img[1155]), .QB(n31336) );
  DFFS img_reg_4__15__3_ ( .D(n12121), .CK(clk), .Q(img[1411]), .QB(n31352) );
  DFFS img_reg_1__15__3_ ( .D(n11735), .CK(clk), .Q(img[1795]), .QB(n31362) );
  DFFS img_reg_13__12__6_ ( .D(n13246), .CK(clk), .Q(img[286]), .QB(n30424) );
  DFFS img_reg_13__10__1_ ( .D(n13235), .CK(clk), .Q(img[297]), .QB(n31135) );
  DFFS img_reg_13__5__1_ ( .D(n13189), .CK(clk), .Q(img[337]), .QB(n31136) );
  DFFS img_reg_13__3__6_ ( .D(n13178), .CK(clk), .Q(img[358]), .QB(n30423) );
  DFFS img_reg_1__14__1_ ( .D(n11731), .CK(clk), .Q(img[1801]), .QB(n31148) );
  DFFS img_reg_15__10__3_ ( .D(n13489), .CK(clk), .Q(img[43]), .QB(n31319) );
  DFFS img_reg_13__13__3_ ( .D(n13255), .CK(clk), .Q(img[275]), .QB(n31275) );
  DFFS img_reg_8__8__3_ ( .D(n12575), .CK(clk), .Q(img[955]), .QB(n31344) );
  DFFS img_reg_4__8__3_ ( .D(n12063), .CK(clk), .Q(img[1467]), .QB(n31354) );
  DFFS img_reg_15__13__3_ ( .D(n13511), .CK(clk), .Q(img[19]), .QB(n31261) );
  DFFS img_reg_5__8__3_ ( .D(n12193), .CK(clk), .Q(img[1339]), .QB(n31342) );
  DFFS img_reg_9__14__3_ ( .D(n12753), .CK(clk), .Q(img[779]), .QB(n31412) );
  DFFS img_reg_13__11__3_ ( .D(n13239), .CK(clk), .Q(img[291]), .QB(n31462) );
  DFFS img_reg_13__10__3_ ( .D(n13233), .CK(clk), .Q(img[299]), .QB(n31325) );
  DFFS img_reg_13__8__3_ ( .D(n13217), .CK(clk), .Q(img[315]), .QB(n31348) );
  DFFS img_reg_13__7__3_ ( .D(n13207), .CK(clk), .Q(img[323]), .QB(n31349) );
  DFFS img_reg_13__6__3_ ( .D(n13201), .CK(clk), .Q(img[331]), .QB(n31426) );
  DFFS img_reg_13__5__3_ ( .D(n13191), .CK(clk), .Q(img[339]), .QB(n31324) );
  DFFS img_reg_13__4__3_ ( .D(n13185), .CK(clk), .Q(img[347]), .QB(n31463) );
  DFFS img_reg_13__3__3_ ( .D(n13175), .CK(clk), .Q(img[355]), .QB(n31490) );
  DFFS img_reg_13__2__3_ ( .D(n13169), .CK(clk), .Q(img[363]), .QB(n31274) );
  DFFS img_reg_13__0__3_ ( .D(n13153), .CK(clk), .Q(img[379]), .QB(n31477) );
  DFFS img_reg_10__13__3_ ( .D(n12873), .CK(clk), .Q(img[659]), .QB(n31284) );
  DFFS img_reg_9__13__3_ ( .D(n12743), .CK(clk), .Q(img[787]), .QB(n31282) );
  DFFS img_reg_8__13__3_ ( .D(n12617), .CK(clk), .Q(img[915]), .QB(n31271) );
  DFFS img_reg_3__14__3_ ( .D(n11985), .CK(clk), .Q(img[1547]), .QB(n31299) );
  DFFS img_reg_12__13__3_ ( .D(n13129), .CK(clk), .Q(img[403]), .QB(n31277) );
  DFFS img_reg_11__13__3_ ( .D(n12999), .CK(clk), .Q(img[531]), .QB(n31259) );
  DFFS img_reg_13__9__3_ ( .D(n13223), .CK(clk), .Q(img[307]), .QB(n31425) );
  DFFS img_reg_12__8__7_ ( .D(n13085), .CK(clk), .Q(img[447]), .QB(n30182) );
  DFFS img_reg_15__8__7_ ( .D(n13469), .CK(clk), .Q(img[63]), .QB(n30166) );
  DFFS img_reg_15__7__7_ ( .D(n13467), .CK(clk), .Q(img[71]), .QB(n30167) );
  DFFS img_reg_8__7__7_ ( .D(n12565), .CK(clk), .Q(img[967]), .QB(n30177) );
  DFFS img_reg_6__15__7_ ( .D(n12373), .CK(clk), .Q(img[1159]), .QB(n30168) );
  DFFS img_reg_5__15__7_ ( .D(n12251), .CK(clk), .Q(img[1287]), .QB(n30172) );
  DFFS img_reg_4__15__7_ ( .D(n12117), .CK(clk), .Q(img[1415]), .QB(n30184) );
  DFFS img_reg_4__8__7_ ( .D(n12067), .CK(clk), .Q(img[1471]), .QB(n30186) );
  DFFS img_reg_5__8__7_ ( .D(n12189), .CK(clk), .Q(img[1343]), .QB(n30174) );
  DFFS img_reg_8__10__5_ ( .D(n12595), .CK(clk), .Q(img[941]), .QB(n30925) );
  DFFS img_reg_8__10__4_ ( .D(n12594), .CK(clk), .Q(img[940]), .QB(n31902) );
  DFFS img_reg_8__10__3_ ( .D(n12593), .CK(clk), .Q(img[939]), .QB(n31321) );
  DFFS img_reg_8__10__1_ ( .D(n12591), .CK(clk), .Q(img[937]), .QB(n31131) );
  DFFS img_reg_13__8__7_ ( .D(n13213), .CK(clk), .Q(img[319]), .QB(n30180) );
  DFFS img_reg_13__7__7_ ( .D(n13211), .CK(clk), .Q(img[327]), .QB(n30181) );
  DFFS img_reg_5__10__4_ ( .D(n12208), .CK(clk), .Q(img[1324]), .QB(n31875) );
  DFFS img_reg_4__10__4_ ( .D(n12080), .CK(clk), .Q(img[1452]), .QB(n31887) );
  DFFS img_reg_6__13__4_ ( .D(n12360), .CK(clk), .Q(img[1172]), .QB(n31873) );
  DFFS img_reg_4__13__4_ ( .D(n12104), .CK(clk), .Q(img[1428]), .QB(n31889) );
  DFFS img_reg_13__13__4_ ( .D(n13256), .CK(clk), .Q(img[276]), .QB(n31883) );
  DFFS img_reg_15__13__4_ ( .D(n13512), .CK(clk), .Q(img[20]), .QB(n31869) );
  DFFS img_reg_10__13__4_ ( .D(n12872), .CK(clk), .Q(img[660]), .QB(n31892) );
  DFFS img_reg_9__13__4_ ( .D(n12744), .CK(clk), .Q(img[788]), .QB(n31891) );
  DFFS img_reg_8__13__4_ ( .D(n12616), .CK(clk), .Q(img[916]), .QB(n31879) );
  DFFS img_reg_7__13__2_ ( .D(n12485), .CK(clk), .Q(img[1042]), .QB(n30618) );
  DFFS img_reg_2__13__2_ ( .D(n11850), .CK(clk), .Q(img[1682]), .QB(n30565) );
  DFFS img_reg_1__13__0_ ( .D(n11724), .CK(clk), .Q(img[1808]), .QB(n31606) );
  DFFS img_reg_4__14__2_ ( .D(n12110), .CK(clk), .Q(img[1418]), .QB(n30551) );
  DFFS img_reg_1__9__2_ ( .D(n11686), .CK(clk), .Q(img[1842]), .QB(n30559) );
  DFFS img_reg_12__13__4_ ( .D(n13128), .CK(clk), .Q(img[404]), .QB(n31885) );
  DFFS img_reg_11__13__4_ ( .D(n13000), .CK(clk), .Q(img[532]), .QB(n31867) );
  DFFS img_reg_1__11__0_ ( .D(n11708), .CK(clk), .Q(img[1824]), .QB(n31501) );
  DFFS img_reg_11__15__0_ ( .D(n13020), .CK(clk), .Q(img[512]), .QB(n31560) );
  DFFS img_reg_3__9__2_ ( .D(n11942), .CK(clk), .Q(img[1586]), .QB(n30575) );
  DFFS img_reg_9__9__2_ ( .D(n12710), .CK(clk), .Q(img[818]), .QB(n30709) );
  DFFS img_reg_9__9__0_ ( .D(n12716), .CK(clk), .Q(img[816]), .QB(n31724) );
  DFFS img_reg_8__9__2_ ( .D(n12586), .CK(clk), .Q(img[946]), .QB(n30703) );
  DFFS img_reg_8__9__0_ ( .D(n12588), .CK(clk), .Q(img[944]), .QB(n31716) );
  DFFS img_reg_5__10__2_ ( .D(n12210), .CK(clk), .Q(img[1322]), .QB(n30601) );
  DFFS img_reg_5__10__0_ ( .D(n12212), .CK(clk), .Q(img[1320]), .QB(n31581) );
  DFFS img_reg_9__3__2_ ( .D(n12662), .CK(clk), .Q(img[866]), .QB(n30757) );
  DFFS img_reg_9__10__2_ ( .D(n12722), .CK(clk), .Q(img[810]), .QB(n30615) );
  DFFS img_reg_9__10__0_ ( .D(n12724), .CK(clk), .Q(img[808]), .QB(n31709) );
  DFFS img_reg_8__10__2_ ( .D(n12592), .CK(clk), .Q(img[938]), .QB(n30603) );
  DFFS img_reg_8__10__0_ ( .D(n12596), .CK(clk), .Q(img[936]), .QB(n31703) );
  DFFS img_reg_4__10__2_ ( .D(n12078), .CK(clk), .Q(img[1450]), .QB(n30613) );
  DFFS img_reg_15__15__0_ ( .D(n13532), .CK(clk), .Q(img[0]), .QB(n31562) );
  DFFS img_reg_7__11__2_ ( .D(n12470), .CK(clk), .Q(img[1058]), .QB(n30739) );
  DFFS img_reg_7__11__0_ ( .D(n12476), .CK(clk), .Q(img[1056]), .QB(n31696) );
  DFFS img_reg_3__11__0_ ( .D(n11964), .CK(clk), .Q(img[1568]), .QB(n31539) );
  DFFS img_reg_10__11__2_ ( .D(n12858), .CK(clk), .Q(img[674]), .QB(n30735) );
  DFFS img_reg_10__11__0_ ( .D(n12860), .CK(clk), .Q(img[672]), .QB(n31692) );
  DFFS img_reg_9__11__2_ ( .D(n12726), .CK(clk), .Q(img[802]), .QB(n30734) );
  DFFS img_reg_9__11__0_ ( .D(n12732), .CK(clk), .Q(img[800]), .QB(n31691) );
  DFFS img_reg_4__11__2_ ( .D(n12090), .CK(clk), .Q(img[1442]), .QB(n30732) );
  DFFS img_reg_4__11__0_ ( .D(n12092), .CK(clk), .Q(img[1440]), .QB(n31689) );
  DFFS img_reg_12__9__2_ ( .D(n13098), .CK(clk), .Q(img[434]), .QB(n30707) );
  DFFS img_reg_12__9__0_ ( .D(n13100), .CK(clk), .Q(img[432]), .QB(n31722) );
  DFFS img_reg_12__6__2_ ( .D(n13070), .CK(clk), .Q(img[458]), .QB(n30708) );
  DFFS img_reg_12__6__0_ ( .D(n13076), .CK(clk), .Q(img[456]), .QB(n31723) );
  DFFS img_reg_7__14__2_ ( .D(n12498), .CK(clk), .Q(img[1034]), .QB(n30582) );
  DFFS img_reg_7__14__0_ ( .D(n12500), .CK(clk), .Q(img[1032]), .QB(n31666) );
  DFFS img_reg_2__14__2_ ( .D(n11854), .CK(clk), .Q(img[1674]), .QB(n30570) );
  DFFS img_reg_2__12__0_ ( .D(n11844), .CK(clk), .Q(img[1688]), .QB(n31533) );
  DFFS img_reg_12__11__2_ ( .D(n13114), .CK(clk), .Q(img[418]), .QB(n30728) );
  DFFS img_reg_12__10__0_ ( .D(n13108), .CK(clk), .Q(img[424]), .QB(n31707) );
  DFFS img_reg_12__8__2_ ( .D(n13087), .CK(clk), .Q(img[442]), .QB(n30770) );
  DFFS img_reg_12__8__0_ ( .D(n13092), .CK(clk), .Q(img[440]), .QB(n31527) );
  DFFS img_reg_15__12__2_ ( .D(n13506), .CK(clk), .Q(img[26]), .QB(n30748) );
  DFFS img_reg_15__12__0_ ( .D(n13508), .CK(clk), .Q(img[24]), .QB(n31729) );
  DFFS img_reg_15__11__2_ ( .D(n13494), .CK(clk), .Q(img[34]), .QB(n30714) );
  DFFS img_reg_15__8__2_ ( .D(n13474), .CK(clk), .Q(img[58]), .QB(n30762) );
  DFFS img_reg_15__8__0_ ( .D(n13476), .CK(clk), .Q(img[56]), .QB(n31515) );
  DFFS img_reg_15__7__2_ ( .D(n13462), .CK(clk), .Q(img[66]), .QB(n30763) );
  DFFS img_reg_15__7__0_ ( .D(n13468), .CK(clk), .Q(img[64]), .QB(n31516) );
  DFFS img_reg_15__6__2_ ( .D(n13458), .CK(clk), .Q(img[74]), .QB(n30702) );
  DFFS img_reg_15__6__0_ ( .D(n13460), .CK(clk), .Q(img[72]), .QB(n31715) );
  DFFS img_reg_15__5__2_ ( .D(n13446), .CK(clk), .Q(img[82]), .QB(n30594) );
  DFFS img_reg_15__5__0_ ( .D(n13452), .CK(clk), .Q(img[80]), .QB(n31702) );
  DFFS img_reg_12__12__2_ ( .D(n13118), .CK(clk), .Q(img[410]), .QB(n30756) );
  DFFS img_reg_12__12__0_ ( .D(n13124), .CK(clk), .Q(img[408]), .QB(n31737) );
  DFFS img_reg_7__12__2_ ( .D(n12482), .CK(clk), .Q(img[1050]), .QB(n30737) );
  DFFS img_reg_7__12__0_ ( .D(n12484), .CK(clk), .Q(img[1048]), .QB(n31694) );
  DFFS img_reg_1__12__0_ ( .D(n11716), .CK(clk), .Q(img[1816]), .QB(n31503) );
  DFFS img_reg_15__4__2_ ( .D(n13442), .CK(clk), .Q(img[90]), .QB(n30715) );
  DFFS img_reg_15__3__2_ ( .D(n13430), .CK(clk), .Q(img[98]), .QB(n30747) );
  DFFS img_reg_15__3__0_ ( .D(n13436), .CK(clk), .Q(img[96]), .QB(n31730) );
  DFFS img_reg_15__1__2_ ( .D(n13414), .CK(clk), .Q(img[114]), .QB(n30530) );
  DFFS img_reg_15__0__2_ ( .D(n13410), .CK(clk), .Q(img[122]), .QB(n30696) );
  DFFS img_reg_15__0__0_ ( .D(n13412), .CK(clk), .Q(img[120]), .QB(n31561) );
  DFFS img_reg_15__2__2_ ( .D(n13426), .CK(clk), .Q(img[106]), .QB(n30628) );
  DFFS img_reg_15__2__0_ ( .D(n13428), .CK(clk), .Q(img[104]), .QB(n31576) );
  DFFS img_reg_11__12__2_ ( .D(n12994), .CK(clk), .Q(img[538]), .QB(n30746) );
  DFFS img_reg_11__12__0_ ( .D(n12996), .CK(clk), .Q(img[536]), .QB(n31727) );
  DFFS img_reg_10__12__2_ ( .D(n12862), .CK(clk), .Q(img[666]), .QB(n30760) );
  DFFS img_reg_10__12__0_ ( .D(n12868), .CK(clk), .Q(img[664]), .QB(n31740) );
  DFFS img_reg_9__12__2_ ( .D(n12738), .CK(clk), .Q(img[794]), .QB(n30758) );
  DFFS img_reg_9__12__0_ ( .D(n12740), .CK(clk), .Q(img[792]), .QB(n31739) );
  DFFS img_reg_8__12__2_ ( .D(n12606), .CK(clk), .Q(img[922]), .QB(n30750) );
  DFFS img_reg_8__12__0_ ( .D(n12612), .CK(clk), .Q(img[920]), .QB(n31731) );
  DFFS img_reg_6__12__2_ ( .D(n12350), .CK(clk), .Q(img[1178]), .QB(n30716) );
  DFFS img_reg_6__12__0_ ( .D(n12356), .CK(clk), .Q(img[1176]), .QB(n31671) );
  DFFS img_reg_6__10__2_ ( .D(n12334), .CK(clk), .Q(img[1194]), .QB(n30597) );
  DFFS img_reg_6__10__0_ ( .D(n12340), .CK(clk), .Q(img[1192]), .QB(n31577) );
  DFFS img_reg_8__7__2_ ( .D(n12570), .CK(clk), .Q(img[962]), .QB(n30765) );
  DFFS img_reg_8__7__0_ ( .D(n12572), .CK(clk), .Q(img[960]), .QB(n31522) );
  DFFS img_reg_8__6__2_ ( .D(n12558), .CK(clk), .Q(img[970]), .QB(n30704) );
  DFFS img_reg_8__6__0_ ( .D(n12564), .CK(clk), .Q(img[968]), .QB(n31717) );
  DFFS img_reg_8__5__2_ ( .D(n12554), .CK(clk), .Q(img[978]), .QB(n30604) );
  DFFS img_reg_8__5__0_ ( .D(n12556), .CK(clk), .Q(img[976]), .QB(n31704) );
  DFFS img_reg_8__4__2_ ( .D(n12542), .CK(clk), .Q(img[986]), .QB(n30744) );
  DFFS img_reg_8__4__0_ ( .D(n12548), .CK(clk), .Q(img[984]), .QB(n31680) );
  DFFS img_reg_8__3__2_ ( .D(n12538), .CK(clk), .Q(img[994]), .QB(n30749) );
  DFFS img_reg_8__3__0_ ( .D(n12540), .CK(clk), .Q(img[992]), .QB(n31732) );
  DFFS img_reg_8__2__2_ ( .D(n12526), .CK(clk), .Q(img[1002]), .QB(n30630) );
  DFFS img_reg_8__2__0_ ( .D(n12532), .CK(clk), .Q(img[1000]), .QB(n31586) );
  DFFS img_reg_8__1__2_ ( .D(n12522), .CK(clk), .Q(img[1010]), .QB(n30540) );
  DFFS img_reg_8__1__0_ ( .D(n12524), .CK(clk), .Q(img[1008]), .QB(n31648) );
  DFFS img_reg_8__0__2_ ( .D(n12510), .CK(clk), .Q(img[1018]), .QB(n30698) );
  DFFS img_reg_8__0__0_ ( .D(n12516), .CK(clk), .Q(img[1016]), .QB(n31563) );
  DFFS img_reg_6__13__2_ ( .D(n12362), .CK(clk), .Q(img[1170]), .QB(n30595) );
  DFFS img_reg_6__13__0_ ( .D(n12364), .CK(clk), .Q(img[1168]), .QB(n31579) );
  DFFS img_reg_4__13__2_ ( .D(n12106), .CK(clk), .Q(img[1426]), .QB(n30611) );
  DFFS img_reg_4__13__0_ ( .D(n12108), .CK(clk), .Q(img[1424]), .QB(n31595) );
  DFFS img_reg_13__15__0_ ( .D(n13276), .CK(clk), .Q(img[256]), .QB(n31568) );
  DFFS img_reg_10__15__0_ ( .D(n12892), .CK(clk), .Q(img[640]), .QB(n31572) );
  DFFS img_reg_9__15__0_ ( .D(n12764), .CK(clk), .Q(img[768]), .QB(n31570) );
  DFFS img_reg_8__15__0_ ( .D(n12636), .CK(clk), .Q(img[896]), .QB(n31564) );
  DFFS img_reg_6__15__2_ ( .D(n12378), .CK(clk), .Q(img[1154]), .QB(n30639) );
  DFFS img_reg_6__15__0_ ( .D(n12380), .CK(clk), .Q(img[1152]), .QB(n31497) );
  DFFS img_reg_5__15__0_ ( .D(n12252), .CK(clk), .Q(img[1280]), .QB(n31517) );
  DFFS img_reg_4__15__0_ ( .D(n12124), .CK(clk), .Q(img[1408]), .QB(n31511) );
  DFFS img_reg_3__15__0_ ( .D(n11996), .CK(clk), .Q(img[1536]), .QB(n31543) );
  DFFS img_reg_2__15__0_ ( .D(n11868), .CK(clk), .Q(img[1664]), .QB(n31535) );
  DFFS img_reg_1__15__0_ ( .D(n11740), .CK(clk), .Q(img[1792]), .QB(n31505) );
  DFFS img_reg_0__15__0_ ( .D(n11612), .CK(clk), .Q(img[1920]), .QB(n31555) );
  DFFS img_reg_15__10__2_ ( .D(n13490), .CK(clk), .Q(img[42]), .QB(n30593) );
  DFFS img_reg_15__10__0_ ( .D(n13492), .CK(clk), .Q(img[40]), .QB(n31701) );
  DFFS img_reg_6__9__2_ ( .D(n12330), .CK(clk), .Q(img[1202]), .QB(n30532) );
  DFFS img_reg_4__9__2_ ( .D(n12074), .CK(clk), .Q(img[1458]), .QB(n30548) );
  DFFS img_reg_13__13__2_ ( .D(n13254), .CK(clk), .Q(img[274]), .QB(n30625) );
  DFFS img_reg_13__13__0_ ( .D(n13260), .CK(clk), .Q(img[272]), .QB(n31589) );
  DFFS img_reg_8__8__0_ ( .D(n12580), .CK(clk), .Q(img[952]), .QB(n31521) );
  DFFS img_reg_4__8__0_ ( .D(n12068), .CK(clk), .Q(img[1464]), .QB(n31513) );
  DFFS img_reg_15__13__2_ ( .D(n13510), .CK(clk), .Q(img[18]), .QB(n30629) );
  DFFS img_reg_15__13__0_ ( .D(n13516), .CK(clk), .Q(img[16]), .QB(n31575) );
  DFFS img_reg_7__8__0_ ( .D(n12452), .CK(clk), .Q(img[1080]), .QB(n31549) );
  DFFS img_reg_5__8__0_ ( .D(n12196), .CK(clk), .Q(img[1336]), .QB(n31519) );
  DFFS img_reg_3__8__0_ ( .D(n11940), .CK(clk), .Q(img[1592]), .QB(n31545) );
  DFFS img_reg_2__8__0_ ( .D(n11812), .CK(clk), .Q(img[1720]), .QB(n31537) );
  DFFS img_reg_15__9__2_ ( .D(n13483), .CK(clk), .Q(img[50]), .QB(n30701) );
  DFFS img_reg_15__9__0_ ( .D(n13484), .CK(clk), .Q(img[48]), .QB(n31714) );
  DFFS img_reg_11__14__2_ ( .D(n13010), .CK(clk), .Q(img[522]), .QB(n30529) );
  DFFS img_reg_10__14__2_ ( .D(n12878), .CK(clk), .Q(img[650]), .QB(n30554) );
  DFFS img_reg_10__14__0_ ( .D(n12884), .CK(clk), .Q(img[648]), .QB(n31662) );
  DFFS img_reg_9__14__2_ ( .D(n12754), .CK(clk), .Q(img[778]), .QB(n30552) );
  DFFS img_reg_6__14__2_ ( .D(n12366), .CK(clk), .Q(img[1162]), .QB(n30535) );
  DFFS img_reg_13__12__2_ ( .D(n13250), .CK(clk), .Q(img[282]), .QB(n30754) );
  DFFS img_reg_13__12__0_ ( .D(n13252), .CK(clk), .Q(img[280]), .QB(n31735) );
  DFFS img_reg_13__11__2_ ( .D(n13238), .CK(clk), .Q(img[290]), .QB(n30726) );
  DFFS img_reg_13__11__0_ ( .D(n13244), .CK(clk), .Q(img[288]), .QB(n31683) );
  DFFS img_reg_13__10__2_ ( .D(n13234), .CK(clk), .Q(img[298]), .QB(n30607) );
  DFFS img_reg_13__10__0_ ( .D(n13236), .CK(clk), .Q(img[296]), .QB(n31705) );
  DFFS img_reg_13__8__2_ ( .D(n13218), .CK(clk), .Q(img[314]), .QB(n30768) );
  DFFS img_reg_13__8__0_ ( .D(n13220), .CK(clk), .Q(img[312]), .QB(n31525) );
  DFFS img_reg_13__7__2_ ( .D(n13206), .CK(clk), .Q(img[322]), .QB(n30769) );
  DFFS img_reg_13__7__0_ ( .D(n13212), .CK(clk), .Q(img[320]), .QB(n31526) );
  DFFS img_reg_13__6__2_ ( .D(n13202), .CK(clk), .Q(img[330]), .QB(n30711) );
  DFFS img_reg_13__6__0_ ( .D(n13204), .CK(clk), .Q(img[328]), .QB(n31721) );
  DFFS img_reg_13__5__2_ ( .D(n13190), .CK(clk), .Q(img[338]), .QB(n30608) );
  DFFS img_reg_13__4__2_ ( .D(n13186), .CK(clk), .Q(img[346]), .QB(n30727) );
  DFFS img_reg_13__4__0_ ( .D(n13188), .CK(clk), .Q(img[344]), .QB(n31684) );
  DFFS img_reg_13__3__2_ ( .D(n13174), .CK(clk), .Q(img[354]), .QB(n30753) );
  DFFS img_reg_13__3__0_ ( .D(n13180), .CK(clk), .Q(img[352]), .QB(n31736) );
  DFFS img_reg_13__2__2_ ( .D(n13170), .CK(clk), .Q(img[362]), .QB(n30624) );
  DFFS img_reg_13__2__0_ ( .D(n13172), .CK(clk), .Q(img[360]), .QB(n31590) );
  DFFS img_reg_13__1__2_ ( .D(n13158), .CK(clk), .Q(img[370]), .QB(n30544) );
  DFFS img_reg_13__0__0_ ( .D(n13156), .CK(clk), .Q(img[376]), .QB(n31567) );
  DFFS img_reg_10__13__2_ ( .D(n12874), .CK(clk), .Q(img[658]), .QB(n30623) );
  DFFS img_reg_10__13__0_ ( .D(n12876), .CK(clk), .Q(img[656]), .QB(n31598) );
  DFFS img_reg_9__13__2_ ( .D(n12742), .CK(clk), .Q(img[786]), .QB(n30636) );
  DFFS img_reg_9__13__0_ ( .D(n12748), .CK(clk), .Q(img[784]), .QB(n31597) );
  DFFS img_reg_8__13__2_ ( .D(n12618), .CK(clk), .Q(img[914]), .QB(n30631) );
  DFFS img_reg_8__13__0_ ( .D(n12620), .CK(clk), .Q(img[912]), .QB(n31585) );
  DFFS img_reg_5__14__2_ ( .D(n12242), .CK(clk), .Q(img[1290]), .QB(n30539) );
  DFFS img_reg_3__14__2_ ( .D(n11986), .CK(clk), .Q(img[1546]), .QB(n30578) );
  DFFS img_reg_1__14__2_ ( .D(n11730), .CK(clk), .Q(img[1802]), .QB(n30562) );
  DFFS img_reg_1__14__0_ ( .D(n11732), .CK(clk), .Q(img[1800]), .QB(n31602) );
  DFFS img_reg_12__13__2_ ( .D(n13130), .CK(clk), .Q(img[402]), .QB(n30635) );
  DFFS img_reg_12__13__0_ ( .D(n13132), .CK(clk), .Q(img[400]), .QB(n31591) );
  DFFS img_reg_11__13__2_ ( .D(n12998), .CK(clk), .Q(img[530]), .QB(n30627) );
  DFFS img_reg_11__13__0_ ( .D(n13004), .CK(clk), .Q(img[528]), .QB(n31573) );
  DFFS img_reg_13__9__2_ ( .D(n13222), .CK(clk), .Q(img[306]), .QB(n30710) );
  DFFS img_reg_13__9__0_ ( .D(n13228), .CK(clk), .Q(img[304]), .QB(n31720) );
  DFFS img_reg_10__10__5_ ( .D(n12849), .CK(clk), .Q(img[685]), .QB(n30935) );
  DFFS img_reg_10__10__3_ ( .D(n12847), .CK(clk), .Q(img[683]), .QB(n31331) );
  DFFS img_reg_10__10__2_ ( .D(n12846), .CK(clk), .Q(img[682]), .QB(n30616) );
  DFFS img_reg_10__10__1_ ( .D(n12845), .CK(clk), .Q(img[681]), .QB(n31144) );
  DFFS img_reg_8__11__6_ ( .D(n12598), .CK(clk), .Q(img[934]), .QB(n30457) );
  DFFS img_reg_8__11__5_ ( .D(n12599), .CK(clk), .Q(img[933]), .QB(n30999) );
  DFFS img_reg_8__11__3_ ( .D(n12601), .CK(clk), .Q(img[931]), .QB(n31452) );
  DFFS img_reg_8__11__2_ ( .D(n12602), .CK(clk), .Q(img[930]), .QB(n30743) );
  DFFS img_reg_8__11__0_ ( .D(n12604), .CK(clk), .Q(img[928]), .QB(n31679) );
  DFFS img_reg_0__9__5_ ( .D(n11559), .CK(clk), .Q(img[1973]), .QB(n30887) );
  DFFS img_reg_0__9__3_ ( .D(n11561), .CK(clk), .Q(img[1971]), .QB(n31309) );
  DFFS img_reg_0__9__2_ ( .D(n11562), .CK(clk), .Q(img[1970]), .QB(n30587) );
  DFFS img_reg_0__9__1_ ( .D(n11563), .CK(clk), .Q(img[1969]), .QB(n31174) );
  DFFS img_reg_0__9__0_ ( .D(n11564), .CK(clk), .Q(img[1968]), .QB(n31628) );
  DFFS img_reg_0__10__5_ ( .D(n11569), .CK(clk), .Q(img[1965]), .QB(n30890) );
  DFFS img_reg_0__10__3_ ( .D(n11567), .CK(clk), .Q(img[1963]), .QB(n31313) );
  DFFS img_reg_0__10__2_ ( .D(n11566), .CK(clk), .Q(img[1962]), .QB(n30583) );
  DFFS img_reg_0__10__0_ ( .D(n11572), .CK(clk), .Q(img[1960]), .QB(n31632) );
  DFFS img_reg_7__13__6_ ( .D(n12489), .CK(clk), .Q(img[1046]), .QB(n30490) );
  DFFS img_reg_2__13__6_ ( .D(n11846), .CK(clk), .Q(img[1686]), .QB(n30381) );
  DFFS img_reg_2__13__1_ ( .D(n11851), .CK(clk), .Q(img[1681]), .QB(n31158) );
  DFFS img_reg_7__9__6_ ( .D(n12458), .CK(clk), .Q(img[1078]), .QB(n30395) );
  DFFS img_reg_7__9__1_ ( .D(n12453), .CK(clk), .Q(img[1073]), .QB(n31207) );
  DFFS img_reg_1__9__6_ ( .D(n11690), .CK(clk), .Q(img[1846]), .QB(n30375) );
  DFFS img_reg_1__11__6_ ( .D(n11706), .CK(clk), .Q(img[1830]), .QB(n30308) );
  DFFS img_reg_1__11__1_ ( .D(n11701), .CK(clk), .Q(img[1825]), .QB(n31038) );
  DFFS img_reg_2__10__5_ ( .D(n11825), .CK(clk), .Q(img[1709]), .QB(n30871) );
  DFFS img_reg_2__10__3_ ( .D(n11823), .CK(clk), .Q(img[1707]), .QB(n31293) );
  DFFS img_reg_2__10__2_ ( .D(n11822), .CK(clk), .Q(img[1706]), .QB(n30563) );
  DFFS img_reg_2__10__1_ ( .D(n11821), .CK(clk), .Q(img[1705]), .QB(n31160) );
  DFFS img_reg_2__10__0_ ( .D(n11828), .CK(clk), .Q(img[1704]), .QB(n31612) );
  DFFS img_reg_12__15__6_ ( .D(n13142), .CK(clk), .Q(img[390]), .QB(n30468) );
  DFFS img_reg_12__15__1_ ( .D(n13147), .CK(clk), .Q(img[385]), .QB(n31029) );
  DFFS img_reg_11__15__6_ ( .D(n13018), .CK(clk), .Q(img[518]), .QB(n30471) );
  DFFS img_reg_11__15__1_ ( .D(n13013), .CK(clk), .Q(img[513]), .QB(n31012) );
  DFFS img_reg_3__9__6_ ( .D(n11946), .CK(clk), .Q(img[1590]), .QB(n30391) );
  DFFS img_reg_8__9__1_ ( .D(n12587), .CK(clk), .Q(img[945]), .QB(n31217) );
  DFFS img_reg_5__10__6_ ( .D(n12206), .CK(clk), .Q(img[1326]), .QB(n30485) );
  DFFS img_reg_0__9__6_ ( .D(n11558), .CK(clk), .Q(img[1974]), .QB(n30403) );
  DFFS img_reg_9__6__1_ ( .D(n12691), .CK(clk), .Q(img[841]), .QB(n31226) );
  DFFS img_reg_9__0__1_ ( .D(n12643), .CK(clk), .Q(img[889]), .QB(n31034) );
  DFFS img_reg_10__10__6_ ( .D(n12850), .CK(clk), .Q(img[686]), .QB(n30512) );
  DFFS img_reg_9__10__6_ ( .D(n12718), .CK(clk), .Q(img[814]), .QB(n30510) );
  DFFS img_reg_8__10__6_ ( .D(n12590), .CK(clk), .Q(img[942]), .QB(n30503) );
  DFFS img_reg_4__10__6_ ( .D(n12082), .CK(clk), .Q(img[1454]), .QB(n30489) );
  DFFS img_reg_15__15__6_ ( .D(n13526), .CK(clk), .Q(img[6]), .QB(n30473) );
  DFFS img_reg_15__15__1_ ( .D(n13531), .CK(clk), .Q(img[1]), .QB(n31014) );
  DFFS img_reg_2__10__6_ ( .D(n11826), .CK(clk), .Q(img[1710]), .QB(n30379) );
  DFFS img_reg_0__10__6_ ( .D(n11570), .CK(clk), .Q(img[1966]), .QB(n30399) );
  DFFS img_reg_7__11__6_ ( .D(n12474), .CK(clk), .Q(img[1062]), .QB(n30434) );
  DFFS img_reg_3__11__6_ ( .D(n11962), .CK(clk), .Q(img[1574]), .QB(n30324) );
  DFFS img_reg_3__11__1_ ( .D(n11957), .CK(clk), .Q(img[1569]), .QB(n31054) );
  DFFS img_reg_10__11__6_ ( .D(n12854), .CK(clk), .Q(img[678]), .QB(n30466) );
  DFFS img_reg_10__11__1_ ( .D(n12859), .CK(clk), .Q(img[673]), .QB(n31099) );
  DFFS img_reg_9__11__6_ ( .D(n12730), .CK(clk), .Q(img[806]), .QB(n30465) );
  DFFS img_reg_9__11__1_ ( .D(n12725), .CK(clk), .Q(img[801]), .QB(n31097) );
  DFFS img_reg_8__11__1_ ( .D(n12603), .CK(clk), .Q(img[929]), .QB(n31086) );
  DFFS img_reg_4__11__1_ ( .D(n12091), .CK(clk), .Q(img[1441]), .QB(n31096) );
  DFFS img_reg_12__9__6_ ( .D(n13094), .CK(clk), .Q(img[438]), .QB(n30448) );
  DFFS img_reg_12__9__1_ ( .D(n13099), .CK(clk), .Q(img[433]), .QB(n31223) );
  DFFS img_reg_12__6__6_ ( .D(n13074), .CK(clk), .Q(img[462]), .QB(n30449) );
  DFFS img_reg_12__6__1_ ( .D(n13069), .CK(clk), .Q(img[457]), .QB(n31224) );
  DFFS img_reg_15__14__6_ ( .D(n13518), .CK(clk), .Q(img[14]), .QB(n30346) );
  DFFS img_reg_7__14__6_ ( .D(n12494), .CK(clk), .Q(img[1038]), .QB(n30397) );
  DFFS img_reg_7__14__1_ ( .D(n12499), .CK(clk), .Q(img[1033]), .QB(n31209) );
  DFFS img_reg_2__14__6_ ( .D(n11858), .CK(clk), .Q(img[1678]), .QB(n30385) );
  DFFS img_reg_2__12__6_ ( .D(n11842), .CK(clk), .Q(img[1694]), .QB(n30318) );
  DFFS img_reg_2__12__1_ ( .D(n11837), .CK(clk), .Q(img[1689]), .QB(n31048) );
  DFFS img_reg_14__13__6_ ( .D(n13382), .CK(clk), .Q(img[150]), .QB(n30519) );
  DFFS img_reg_12__8__6_ ( .D(n13091), .CK(clk), .Q(img[446]), .QB(n30300) );
  DFFS img_reg_12__8__1_ ( .D(n13086), .CK(clk), .Q(img[441]), .QB(n31240) );
  DFFS img_reg_15__12__1_ ( .D(n13507), .CK(clk), .Q(img[25]), .QB(n31107) );
  DFFS img_reg_15__11__6_ ( .D(n13498), .CK(clk), .Q(img[38]), .QB(n30455) );
  DFFS img_reg_15__11__1_ ( .D(n13493), .CK(clk), .Q(img[33]), .QB(n31076) );
  DFFS img_reg_15__8__6_ ( .D(n13470), .CK(clk), .Q(img[62]), .QB(n30284) );
  DFFS img_reg_15__8__1_ ( .D(n13475), .CK(clk), .Q(img[57]), .QB(n31232) );
  DFFS img_reg_15__7__6_ ( .D(n13466), .CK(clk), .Q(img[70]), .QB(n30285) );
  DFFS img_reg_15__7__1_ ( .D(n13461), .CK(clk), .Q(img[65]), .QB(n31231) );
  DFFS img_reg_15__6__6_ ( .D(n13454), .CK(clk), .Q(img[78]), .QB(n30441) );
  DFFS img_reg_15__6__1_ ( .D(n13459), .CK(clk), .Q(img[73]), .QB(n31216) );
  DFFS img_reg_15__5__6_ ( .D(n13450), .CK(clk), .Q(img[86]), .QB(n30496) );
  DFFS img_reg_15__5__1_ ( .D(n13445), .CK(clk), .Q(img[81]), .QB(n31122) );
  DFFS img_reg_12__12__1_ ( .D(n13117), .CK(clk), .Q(img[409]), .QB(n31115) );
  DFFS img_reg_7__12__1_ ( .D(n12483), .CK(clk), .Q(img[1049]), .QB(n31100) );
  DFFS img_reg_3__12__6_ ( .D(n11966), .CK(clk), .Q(img[1566]), .QB(n30326) );
  DFFS img_reg_3__12__1_ ( .D(n11971), .CK(clk), .Q(img[1561]), .QB(n31056) );
  DFFS img_reg_1__12__6_ ( .D(n11710), .CK(clk), .Q(img[1822]), .QB(n30310) );
  DFFS img_reg_1__12__1_ ( .D(n11715), .CK(clk), .Q(img[1817]), .QB(n31040) );
  DFFS img_reg_15__4__1_ ( .D(n13443), .CK(clk), .Q(img[89]), .QB(n31075) );
  DFFS img_reg_15__3__1_ ( .D(n13429), .CK(clk), .Q(img[97]), .QB(n31106) );
  DFFS img_reg_15__1__6_ ( .D(n13418), .CK(clk), .Q(img[118]), .QB(n30347) );
  DFFS img_reg_15__0__6_ ( .D(n13406), .CK(clk), .Q(img[126]), .QB(n30474) );
  DFFS img_reg_15__0__1_ ( .D(n13411), .CK(clk), .Q(img[121]), .QB(n31013) );
  DFFS img_reg_15__2__6_ ( .D(n13422), .CK(clk), .Q(img[110]), .QB(n30516) );
  DFFS img_reg_15__2__1_ ( .D(n13427), .CK(clk), .Q(img[105]), .QB(n31245) );
  DFFS img_reg_11__12__1_ ( .D(n12995), .CK(clk), .Q(img[537]), .QB(n31105) );
  DFFS img_reg_10__12__1_ ( .D(n12861), .CK(clk), .Q(img[665]), .QB(n31118) );
  DFFS img_reg_9__12__1_ ( .D(n12739), .CK(clk), .Q(img[793]), .QB(n31116) );
  DFFS img_reg_8__12__1_ ( .D(n12605), .CK(clk), .Q(img[921]), .QB(n31109) );
  DFFS img_reg_6__12__1_ ( .D(n12349), .CK(clk), .Q(img[1177]), .QB(n31077) );
  DFFS img_reg_6__10__6_ ( .D(n12338), .CK(clk), .Q(img[1198]), .QB(n30501) );
  DFFS img_reg_6__10__1_ ( .D(n12333), .CK(clk), .Q(img[1193]), .QB(n31125) );
  DFFS img_reg_8__7__6_ ( .D(n12566), .CK(clk), .Q(img[966]), .QB(n30295) );
  DFFS img_reg_8__7__1_ ( .D(n12571), .CK(clk), .Q(img[961]), .QB(n31233) );
  DFFS img_reg_8__6__1_ ( .D(n12557), .CK(clk), .Q(img[969]), .QB(n31218) );
  DFFS img_reg_8__5__6_ ( .D(n12550), .CK(clk), .Q(img[982]), .QB(n30502) );
  DFFS img_reg_8__4__6_ ( .D(n12546), .CK(clk), .Q(img[990]), .QB(n30458) );
  DFFS img_reg_8__4__1_ ( .D(n12541), .CK(clk), .Q(img[985]), .QB(n31085) );
  DFFS img_reg_8__3__1_ ( .D(n12539), .CK(clk), .Q(img[993]), .QB(n31108) );
  DFFS img_reg_8__2__6_ ( .D(n12530), .CK(clk), .Q(img[1006]), .QB(n30518) );
  DFFS img_reg_8__2__1_ ( .D(n12525), .CK(clk), .Q(img[1001]), .QB(n31247) );
  DFFS img_reg_8__1__6_ ( .D(n12518), .CK(clk), .Q(img[1014]), .QB(n30357) );
  DFFS img_reg_8__1__1_ ( .D(n12523), .CK(clk), .Q(img[1009]), .QB(n31212) );
  DFFS img_reg_8__0__6_ ( .D(n12514), .CK(clk), .Q(img[1022]), .QB(n30476) );
  DFFS img_reg_8__0__1_ ( .D(n12509), .CK(clk), .Q(img[1017]), .QB(n31023) );
  DFFS img_reg_6__13__6_ ( .D(n12358), .CK(clk), .Q(img[1174]), .QB(n30498) );
  DFFS img_reg_6__13__1_ ( .D(n12363), .CK(clk), .Q(img[1169]), .QB(n31123) );
  DFFS img_reg_4__13__6_ ( .D(n12102), .CK(clk), .Q(img[1430]), .QB(n30486) );
  DFFS img_reg_13__15__6_ ( .D(n13274), .CK(clk), .Q(img[262]), .QB(n30469) );
  DFFS img_reg_13__15__1_ ( .D(n13269), .CK(clk), .Q(img[257]), .QB(n31028) );
  DFFS img_reg_10__15__6_ ( .D(n12886), .CK(clk), .Q(img[646]), .QB(n30480) );
  DFFS img_reg_10__15__1_ ( .D(n12891), .CK(clk), .Q(img[641]), .QB(n31037) );
  DFFS img_reg_9__15__6_ ( .D(n12762), .CK(clk), .Q(img[774]), .QB(n30479) );
  DFFS img_reg_8__15__6_ ( .D(n12630), .CK(clk), .Q(img[902]), .QB(n30475) );
  DFFS img_reg_8__15__1_ ( .D(n12635), .CK(clk), .Q(img[897]), .QB(n31024) );
  DFFS img_reg_7__15__6_ ( .D(n12506), .CK(clk), .Q(img[1030]), .QB(n30332) );
  DFFS img_reg_7__15__1_ ( .D(n12501), .CK(clk), .Q(img[1025]), .QB(n31065) );
  DFFS img_reg_6__15__6_ ( .D(n12374), .CK(clk), .Q(img[1158]), .QB(n30286) );
  DFFS img_reg_6__15__1_ ( .D(n12379), .CK(clk), .Q(img[1153]), .QB(n31018) );
  DFFS img_reg_5__15__6_ ( .D(n12250), .CK(clk), .Q(img[1286]), .QB(n30290) );
  DFFS img_reg_5__15__1_ ( .D(n12245), .CK(clk), .Q(img[1281]), .QB(n31022) );
  DFFS img_reg_4__15__6_ ( .D(n12118), .CK(clk), .Q(img[1414]), .QB(n30302) );
  DFFS img_reg_4__15__1_ ( .D(n12123), .CK(clk), .Q(img[1409]), .QB(n31033) );
  DFFS img_reg_3__15__6_ ( .D(n11994), .CK(clk), .Q(img[1542]), .QB(n30328) );
  DFFS img_reg_3__15__1_ ( .D(n11989), .CK(clk), .Q(img[1537]), .QB(n31061) );
  DFFS img_reg_2__15__6_ ( .D(n11862), .CK(clk), .Q(img[1670]), .QB(n30320) );
  DFFS img_reg_2__15__1_ ( .D(n11867), .CK(clk), .Q(img[1665]), .QB(n31053) );
  DFFS img_reg_1__15__1_ ( .D(n11733), .CK(clk), .Q(img[1793]), .QB(n31045) );
  DFFS img_reg_0__15__6_ ( .D(n11606), .CK(clk), .Q(img[1926]), .QB(n30340) );
  DFFS img_reg_0__15__1_ ( .D(n11611), .CK(clk), .Q(img[1921]), .QB(n31073) );
  DFFS img_reg_15__10__6_ ( .D(n13486), .CK(clk), .Q(img[46]), .QB(n30497) );
  DFFS img_reg_15__10__1_ ( .D(n13491), .CK(clk), .Q(img[41]), .QB(n31121) );
  DFFS img_reg_6__9__6_ ( .D(n12326), .CK(clk), .Q(img[1206]), .QB(n30348) );
  DFFS img_reg_6__9__1_ ( .D(n12331), .CK(clk), .Q(img[1201]), .QB(n31182) );
  DFFS img_reg_4__9__6_ ( .D(n12070), .CK(clk), .Q(img[1462]), .QB(n30364) );
  DFFS img_reg_4__9__1_ ( .D(n12075), .CK(clk), .Q(img[1457]), .QB(n31201) );
  DFFS img_reg_13__13__6_ ( .D(n13258), .CK(clk), .Q(img[278]), .QB(n30521) );
  DFFS img_reg_13__13__1_ ( .D(n13253), .CK(clk), .Q(img[273]), .QB(n31252) );
  DFFS img_reg_8__8__6_ ( .D(n12578), .CK(clk), .Q(img[958]), .QB(n30294) );
  DFFS img_reg_8__8__1_ ( .D(n12573), .CK(clk), .Q(img[953]), .QB(n31234) );
  DFFS img_reg_4__8__6_ ( .D(n12066), .CK(clk), .Q(img[1470]), .QB(n30304) );
  DFFS img_reg_4__8__1_ ( .D(n12061), .CK(clk), .Q(img[1465]), .QB(n31030) );
  DFFS img_reg_15__13__6_ ( .D(n13514), .CK(clk), .Q(img[22]), .QB(n30515) );
  DFFS img_reg_15__13__1_ ( .D(n13509), .CK(clk), .Q(img[17]), .QB(n31246) );
  DFFS img_reg_7__8__6_ ( .D(n12446), .CK(clk), .Q(img[1086]), .QB(n30334) );
  DFFS img_reg_7__8__1_ ( .D(n12451), .CK(clk), .Q(img[1081]), .QB(n31062) );
  DFFS img_reg_5__8__6_ ( .D(n12190), .CK(clk), .Q(img[1342]), .QB(n30292) );
  DFFS img_reg_5__8__1_ ( .D(n12195), .CK(clk), .Q(img[1337]), .QB(n31019) );
  DFFS img_reg_3__8__6_ ( .D(n11934), .CK(clk), .Q(img[1598]), .QB(n30330) );
  DFFS img_reg_3__8__1_ ( .D(n11939), .CK(clk), .Q(img[1593]), .QB(n31058) );
  DFFS img_reg_2__8__6_ ( .D(n11810), .CK(clk), .Q(img[1726]), .QB(n30322) );
  DFFS img_reg_7__13__7_ ( .D(n12490), .CK(clk), .Q(img[1047]), .QB(n30224) );
  DFFS img_reg_2__13__7_ ( .D(n11845), .CK(clk), .Q(img[1687]), .QB(n30075) );
  DFFS img_reg_12__14__7_ ( .D(n13139), .CK(clk), .Q(img[399]), .QB(n30263) );
  DFFS img_reg_7__9__7_ ( .D(n12459), .CK(clk), .Q(img[1079]), .QB(n30091) );
  DFFS img_reg_1__9__7_ ( .D(n11691), .CK(clk), .Q(img[1847]), .QB(n30071) );
  DFFS img_reg_15__9__1_ ( .D(n13482), .CK(clk), .Q(img[49]), .QB(n31215) );
  DFFS img_reg_1__11__7_ ( .D(n11707), .CK(clk), .Q(img[1831]), .QB(n30132) );
  DFFS img_reg_11__14__6_ ( .D(n13006), .CK(clk), .Q(img[526]), .QB(n30344) );
  DFFS img_reg_11__14__1_ ( .D(n13011), .CK(clk), .Q(img[521]), .QB(n31187) );
  DFFS img_reg_10__14__6_ ( .D(n12882), .CK(clk), .Q(img[654]), .QB(n30369) );
  DFFS img_reg_9__14__6_ ( .D(n12750), .CK(clk), .Q(img[782]), .QB(n30368) );
  DFFS img_reg_8__14__6_ ( .D(n12626), .CK(clk), .Q(img[910]), .QB(n30356) );
  DFFS img_reg_8__14__1_ ( .D(n12621), .CK(clk), .Q(img[905]), .QB(n31211) );
  DFFS img_reg_6__14__6_ ( .D(n12370), .CK(clk), .Q(img[1166]), .QB(n30350) );
  DFFS img_reg_6__14__1_ ( .D(n12365), .CK(clk), .Q(img[1161]), .QB(n31184) );
  DFFS img_reg_13__12__1_ ( .D(n13251), .CK(clk), .Q(img[281]), .QB(n31113) );
  DFFS img_reg_13__11__6_ ( .D(n13242), .CK(clk), .Q(img[294]), .QB(n30461) );
  DFFS img_reg_13__11__1_ ( .D(n13237), .CK(clk), .Q(img[289]), .QB(n31090) );
  DFFS img_reg_13__10__6_ ( .D(n13230), .CK(clk), .Q(img[302]), .QB(n30507) );
  DFFS img_reg_13__8__6_ ( .D(n13214), .CK(clk), .Q(img[318]), .QB(n30298) );
  DFFS img_reg_13__8__1_ ( .D(n13219), .CK(clk), .Q(img[313]), .QB(n31238) );
  DFFS img_reg_13__7__6_ ( .D(n13210), .CK(clk), .Q(img[326]), .QB(n30299) );
  DFFS img_reg_13__7__1_ ( .D(n13205), .CK(clk), .Q(img[321]), .QB(n31237) );
  DFFS img_reg_13__6__1_ ( .D(n13203), .CK(clk), .Q(img[329]), .QB(n31222) );
  DFFS img_reg_13__4__6_ ( .D(n13182), .CK(clk), .Q(img[350]), .QB(n30462) );
  DFFS img_reg_13__4__1_ ( .D(n13187), .CK(clk), .Q(img[345]), .QB(n31089) );
  DFFS img_reg_13__3__1_ ( .D(n13173), .CK(clk), .Q(img[353]), .QB(n31112) );
  DFFS img_reg_13__2__6_ ( .D(n13166), .CK(clk), .Q(img[366]), .QB(n30522) );
  DFFS img_reg_13__2__1_ ( .D(n13171), .CK(clk), .Q(img[361]), .QB(n31251) );
  DFFS img_reg_13__1__6_ ( .D(n13162), .CK(clk), .Q(img[374]), .QB(n30361) );
  DFFS img_reg_13__1__1_ ( .D(n13157), .CK(clk), .Q(img[369]), .QB(n31198) );
  DFFS img_reg_13__0__6_ ( .D(n13150), .CK(clk), .Q(img[382]), .QB(n30470) );
  DFFS img_reg_13__0__1_ ( .D(n13155), .CK(clk), .Q(img[377]), .QB(n31027) );
  DFFS img_reg_10__13__6_ ( .D(n12870), .CK(clk), .Q(img[662]), .QB(n30526) );
  DFFS img_reg_10__13__1_ ( .D(n12875), .CK(clk), .Q(img[657]), .QB(n31257) );
  DFFS img_reg_9__13__6_ ( .D(n12746), .CK(clk), .Q(img[790]), .QB(n30525) );
  DFFS img_reg_9__13__1_ ( .D(n12741), .CK(clk), .Q(img[785]), .QB(n31255) );
  DFFS img_reg_8__13__6_ ( .D(n12614), .CK(clk), .Q(img[918]), .QB(n30517) );
  DFFS img_reg_14__14__6_ ( .D(n13394), .CK(clk), .Q(img[142]), .QB(n30358) );
  DFFS img_reg_14__14__1_ ( .D(n13389), .CK(clk), .Q(img[137]), .QB(n31195) );
  DFFS img_reg_5__14__6_ ( .D(n12238), .CK(clk), .Q(img[1294]), .QB(n30354) );
  DFFS img_reg_5__14__1_ ( .D(n12243), .CK(clk), .Q(img[1289]), .QB(n31193) );
  DFFS img_reg_3__14__6_ ( .D(n11982), .CK(clk), .Q(img[1550]), .QB(n30393) );
  DFFS img_reg_1__14__6_ ( .D(n11726), .CK(clk), .Q(img[1806]), .QB(n30377) );
  DFFS img_reg_12__15__7_ ( .D(n13141), .CK(clk), .Q(img[391]), .QB(n30278) );
  DFFS img_reg_11__15__7_ ( .D(n13019), .CK(clk), .Q(img[519]), .QB(n30268) );
  DFFS img_reg_3__9__7_ ( .D(n11947), .CK(clk), .Q(img[1591]), .QB(n30087) );
  DFFS img_reg_12__13__6_ ( .D(n13126), .CK(clk), .Q(img[406]), .QB(n30523) );
  DFFS img_reg_12__13__1_ ( .D(n13131), .CK(clk), .Q(img[401]), .QB(n31254) );
  DFFS img_reg_11__13__6_ ( .D(n13002), .CK(clk), .Q(img[534]), .QB(n30513) );
  DFFS img_reg_11__13__1_ ( .D(n12997), .CK(clk), .Q(img[529]), .QB(n31244) );
  DFFS img_reg_13__9__1_ ( .D(n13221), .CK(clk), .Q(img[305]), .QB(n31221) );
  DFFS img_reg_8__9__7_ ( .D(n12581), .CK(clk), .Q(img[951]), .QB(n30050) );
  DFFS img_reg_0__9__7_ ( .D(n11557), .CK(clk), .Q(img[1975]), .QB(n30099) );
  DFFS img_reg_10__10__7_ ( .D(n12851), .CK(clk), .Q(img[687]), .QB(n30237) );
  DFFS img_reg_9__10__7_ ( .D(n12717), .CK(clk), .Q(img[815]), .QB(n30235) );
  DFFS img_reg_8__10__7_ ( .D(n12589), .CK(clk), .Q(img[943]), .QB(n30239) );
  DFFS img_reg_15__15__7_ ( .D(n13525), .CK(clk), .Q(img[7]), .QB(n30270) );
  DFFS img_reg_2__10__7_ ( .D(n11827), .CK(clk), .Q(img[1711]), .QB(n30073) );
  DFFS img_reg_0__10__7_ ( .D(n11571), .CK(clk), .Q(img[1967]), .QB(n30093) );
  DFFS img_reg_7__11__7_ ( .D(n12475), .CK(clk), .Q(img[1063]), .QB(n30152) );
  DFFS img_reg_3__11__7_ ( .D(n11963), .CK(clk), .Q(img[1575]), .QB(n30148) );
  DFFS img_reg_10__11__7_ ( .D(n12853), .CK(clk), .Q(img[679]), .QB(n30253) );
  DFFS img_reg_9__11__7_ ( .D(n12731), .CK(clk), .Q(img[807]), .QB(n30252) );
  DFFS img_reg_8__11__7_ ( .D(n12597), .CK(clk), .Q(img[935]), .QB(n30246) );
  DFFS img_reg_4__11__7_ ( .D(n12085), .CK(clk), .Q(img[1447]), .QB(n30121) );
  DFFS img_reg_12__6__7_ ( .D(n13075), .CK(clk), .Q(img[463]), .QB(n30057) );
  DFFS img_reg_15__14__7_ ( .D(n13517), .CK(clk), .Q(img[15]), .QB(n30282) );
  DFFS img_reg_7__14__7_ ( .D(n12493), .CK(clk), .Q(img[1039]), .QB(n30089) );
  DFFS img_reg_2__14__7_ ( .D(n11859), .CK(clk), .Q(img[1679]), .QB(n30077) );
  DFFS img_reg_15__12__7_ ( .D(n13501), .CK(clk), .Q(img[31]), .QB(n30104) );
  DFFS img_reg_15__6__7_ ( .D(n13453), .CK(clk), .Q(img[79]), .QB(n30041) );
  DFFS img_reg_15__5__7_ ( .D(n13451), .CK(clk), .Q(img[87]), .QB(n30227) );
  DFFS img_reg_7__12__7_ ( .D(n12477), .CK(clk), .Q(img[1055]), .QB(n30155) );
  DFFS img_reg_15__3__7_ ( .D(n13435), .CK(clk), .Q(img[103]), .QB(n30103) );
  DFFS img_reg_15__1__7_ ( .D(n13419), .CK(clk), .Q(img[119]), .QB(n31995) );
  DFFS img_reg_15__0__7_ ( .D(n13405), .CK(clk), .Q(img[127]), .QB(n30271) );
  DFFS img_reg_15__2__7_ ( .D(n13421), .CK(clk), .Q(img[111]), .QB(n30196) );
  DFFS img_reg_11__12__7_ ( .D(n12989), .CK(clk), .Q(img[543]), .QB(n30102) );
  DFFS img_reg_8__12__7_ ( .D(n12611), .CK(clk), .Q(img[927]), .QB(n30114) );
  DFFS img_reg_6__12__7_ ( .D(n12355), .CK(clk), .Q(img[1183]), .QB(n30108) );
  DFFS img_reg_8__6__7_ ( .D(n12563), .CK(clk), .Q(img[975]), .QB(n30051) );
  DFFS img_reg_8__5__7_ ( .D(n12549), .CK(clk), .Q(img[983]), .QB(n30238) );
  DFFS img_reg_8__3__7_ ( .D(n12533), .CK(clk), .Q(img[999]), .QB(n30113) );
  DFFS img_reg_8__0__7_ ( .D(n12515), .CK(clk), .Q(img[1023]), .QB(n30273) );
  DFFS img_reg_13__15__7_ ( .D(n13275), .CK(clk), .Q(img[263]), .QB(n30276) );
  DFFS img_reg_10__15__7_ ( .D(n12885), .CK(clk), .Q(img[647]), .QB(n30280) );
  DFFS img_reg_9__15__7_ ( .D(n12763), .CK(clk), .Q(img[775]), .QB(n30279) );
  DFFS img_reg_8__15__7_ ( .D(n12629), .CK(clk), .Q(img[903]), .QB(n30272) );
  DFFS img_reg_7__15__7_ ( .D(n12507), .CK(clk), .Q(img[1031]), .QB(n30190) );
  DFFS img_reg_3__15__7_ ( .D(n11995), .CK(clk), .Q(img[1543]), .QB(n30146) );
  DFFS img_reg_2__15__7_ ( .D(n11861), .CK(clk), .Q(img[1671]), .QB(n30138) );
  DFFS img_reg_1__15__7_ ( .D(n11739), .CK(clk), .Q(img[1799]), .QB(n30130) );
  DFFS img_reg_15__10__7_ ( .D(n13485), .CK(clk), .Q(img[47]), .QB(n30228) );
  DFFS img_reg_6__9__7_ ( .D(n12325), .CK(clk), .Q(img[1207]), .QB(n30044) );
  DFFS img_reg_4__9__7_ ( .D(n12069), .CK(clk), .Q(img[1463]), .QB(n30060) );
  DFFS img_reg_7__8__7_ ( .D(n12445), .CK(clk), .Q(img[1087]), .QB(n30192) );
  DFFS img_reg_3__8__7_ ( .D(n11933), .CK(clk), .Q(img[1599]), .QB(n30144) );
  DFFS img_reg_2__8__7_ ( .D(n11811), .CK(clk), .Q(img[1727]), .QB(n30136) );
  DFFS img_reg_15__9__7_ ( .D(n13480), .CK(clk), .Q(img[55]), .QB(n30040) );
  DFFS img_reg_11__14__7_ ( .D(n13005), .CK(clk), .Q(img[527]), .QB(n30255) );
  DFFS img_reg_10__14__7_ ( .D(n12883), .CK(clk), .Q(img[655]), .QB(n30266) );
  DFFS img_reg_9__14__7_ ( .D(n12749), .CK(clk), .Q(img[783]), .QB(n30265) );
  DFFS img_reg_8__14__7_ ( .D(n12627), .CK(clk), .Q(img[911]), .QB(n30257) );
  DFFS img_reg_6__14__7_ ( .D(n12371), .CK(clk), .Q(img[1167]), .QB(n30042) );
  DFFS img_reg_13__12__7_ ( .D(n13245), .CK(clk), .Q(img[287]), .QB(n30118) );
  DFFS img_reg_13__11__7_ ( .D(n13243), .CK(clk), .Q(img[295]), .QB(n30240) );
  DFFS img_reg_13__6__7_ ( .D(n13197), .CK(clk), .Q(img[335]), .QB(n30055) );
  DFFS img_reg_13__5__7_ ( .D(n13195), .CK(clk), .Q(img[343]), .QB(n30231) );
  DFFS img_reg_13__4__7_ ( .D(n13181), .CK(clk), .Q(img[351]), .QB(n30241) );
  DFFS img_reg_13__3__7_ ( .D(n13179), .CK(clk), .Q(img[359]), .QB(n30117) );
  DFFS img_reg_13__1__7_ ( .D(n13163), .CK(clk), .Q(img[375]), .QB(n30262) );
  DFFS img_reg_13__0__7_ ( .D(n13149), .CK(clk), .Q(img[383]), .QB(n30277) );
  DFFS img_reg_10__13__7_ ( .D(n12869), .CK(clk), .Q(img[663]), .QB(n30220) );
  DFFS img_reg_9__13__7_ ( .D(n12747), .CK(clk), .Q(img[791]), .QB(n30218) );
  DFFS img_reg_14__14__7_ ( .D(n13395), .CK(clk), .Q(img[143]), .QB(n30259) );
  DFFS img_reg_5__14__7_ ( .D(n12237), .CK(clk), .Q(img[1295]), .QB(n30046) );
  DFFS img_reg_3__14__7_ ( .D(n11981), .CK(clk), .Q(img[1551]), .QB(n30085) );
  DFFS img_reg_1__14__7_ ( .D(n11725), .CK(clk), .Q(img[1807]), .QB(n30069) );
  DFFS img_reg_12__13__7_ ( .D(n13125), .CK(clk), .Q(img[407]), .QB(n30213) );
  DFFS img_reg_13__9__7_ ( .D(n13227), .CK(clk), .Q(img[311]), .QB(n30054) );
  DFFS img_reg_1__11__4_ ( .D(n11704), .CK(clk), .Q(img[1828]), .QB(n31831) );
  DFFS img_reg_12__15__4_ ( .D(n13144), .CK(clk), .Q(img[388]), .QB(n31984) );
  DFFS img_reg_3__9__4_ ( .D(n11944), .CK(clk), .Q(img[1588]), .QB(n31791) );
  DFFS img_reg_9__9__4_ ( .D(n12712), .CK(clk), .Q(img[820]), .QB(n31766) );
  DFFS img_reg_8__9__4_ ( .D(n12584), .CK(clk), .Q(img[948]), .QB(n31754) );
  DFFS img_reg_0__9__4_ ( .D(n11560), .CK(clk), .Q(img[1972]), .QB(n31803) );
  DFFS img_reg_9__3__4_ ( .D(n12664), .CK(clk), .Q(img[868]), .QB(n31928) );
  DFFS img_reg_10__10__4_ ( .D(n12848), .CK(clk), .Q(img[684]), .QB(n31911) );
  DFFS img_reg_15__15__4_ ( .D(n13528), .CK(clk), .Q(img[4]), .QB(n31976) );
  DFFS img_reg_2__10__4_ ( .D(n11824), .CK(clk), .Q(img[1708]), .QB(n31777) );
  DFFS img_reg_0__10__4_ ( .D(n11568), .CK(clk), .Q(img[1964]), .QB(n31797) );
  DFFS img_reg_3__11__4_ ( .D(n11960), .CK(clk), .Q(img[1572]), .QB(n31847) );
  DFFS img_reg_10__11__4_ ( .D(n12856), .CK(clk), .Q(img[676]), .QB(n31973) );
  DFFS img_reg_9__11__4_ ( .D(n12728), .CK(clk), .Q(img[804]), .QB(n31971) );
  DFFS img_reg_8__11__4_ ( .D(n12600), .CK(clk), .Q(img[932]), .QB(n31964) );
  DFFS img_reg_4__11__4_ ( .D(n12088), .CK(clk), .Q(img[1444]), .QB(n31933) );
  DFFS img_reg_12__6__4_ ( .D(n13072), .CK(clk), .Q(img[460]), .QB(n31761) );
  DFFS img_reg_15__14__4_ ( .D(n13520), .CK(clk), .Q(img[12]), .QB(n31947) );
  DFFS img_reg_8__4__4_ ( .D(n12544), .CK(clk), .Q(img[988]), .QB(n31963) );
  DFFS img_reg_8__0__4_ ( .D(n12512), .CK(clk), .Q(img[1020]), .QB(n31979) );
  DFFS img_reg_13__15__4_ ( .D(n13272), .CK(clk), .Q(img[260]), .QB(n31982) );
  DFFS img_reg_10__15__4_ ( .D(n12888), .CK(clk), .Q(img[644]), .QB(n31986) );
  DFFS img_reg_9__15__4_ ( .D(n12760), .CK(clk), .Q(img[772]), .QB(n31985) );
  DFFS img_reg_8__15__4_ ( .D(n12632), .CK(clk), .Q(img[900]), .QB(n31978) );
  DFFS img_reg_7__15__4_ ( .D(n12504), .CK(clk), .Q(img[1028]), .QB(n31855) );
  DFFS img_reg_6__15__4_ ( .D(n12376), .CK(clk), .Q(img[1156]), .QB(n31809) );
  DFFS img_reg_4__15__4_ ( .D(n12120), .CK(clk), .Q(img[1412]), .QB(n31825) );
  DFFS img_reg_3__15__4_ ( .D(n11992), .CK(clk), .Q(img[1540]), .QB(n31851) );
  DFFS img_reg_2__15__4_ ( .D(n11864), .CK(clk), .Q(img[1668]), .QB(n31843) );
  DFFS img_reg_1__15__4_ ( .D(n11736), .CK(clk), .Q(img[1796]), .QB(n31835) );
  DFFS img_reg_0__15__4_ ( .D(n11608), .CK(clk), .Q(img[1924]), .QB(n31863) );
  DFFS img_reg_15__10__4_ ( .D(n13488), .CK(clk), .Q(img[44]), .QB(n31900) );
  DFFS img_reg_6__9__4_ ( .D(n12328), .CK(clk), .Q(img[1204]), .QB(n31748) );
  DFFS img_reg_4__9__4_ ( .D(n12072), .CK(clk), .Q(img[1460]), .QB(n31764) );
  DFFS img_reg_8__8__4_ ( .D(n12576), .CK(clk), .Q(img[956]), .QB(n31818) );
  DFFS img_reg_4__8__4_ ( .D(n12064), .CK(clk), .Q(img[1468]), .QB(n31828) );
  DFFS img_reg_7__8__4_ ( .D(n12448), .CK(clk), .Q(img[1084]), .QB(n31858) );
  DFFS img_reg_5__8__4_ ( .D(n12192), .CK(clk), .Q(img[1340]), .QB(n31816) );
  DFFS img_reg_3__8__4_ ( .D(n11936), .CK(clk), .Q(img[1596]), .QB(n31854) );
  DFFS img_reg_2__8__4_ ( .D(n11808), .CK(clk), .Q(img[1724]), .QB(n31846) );
  DFFS img_reg_11__14__4_ ( .D(n13008), .CK(clk), .Q(img[524]), .QB(n31945) );
  DFFS img_reg_10__14__4_ ( .D(n12880), .CK(clk), .Q(img[652]), .QB(n31958) );
  DFFS img_reg_9__14__4_ ( .D(n12752), .CK(clk), .Q(img[780]), .QB(n31957) );
  DFFS img_reg_8__14__4_ ( .D(n12624), .CK(clk), .Q(img[908]), .QB(n31949) );
  DFFS img_reg_6__14__4_ ( .D(n12368), .CK(clk), .Q(img[1164]), .QB(n31746) );
  DFFS img_reg_13__12__4_ ( .D(n13248), .CK(clk), .Q(img[284]), .QB(n31913) );
  DFFS img_reg_13__11__4_ ( .D(n13240), .CK(clk), .Q(img[292]), .QB(n31968) );
  DFFS img_reg_13__8__4_ ( .D(n13216), .CK(clk), .Q(img[316]), .QB(n31822) );
  DFFS img_reg_13__7__4_ ( .D(n13208), .CK(clk), .Q(img[324]), .QB(n31821) );
  DFFS img_reg_13__6__4_ ( .D(n13200), .CK(clk), .Q(img[332]), .QB(n31759) );
  DFFS img_reg_13__4__4_ ( .D(n13184), .CK(clk), .Q(img[348]), .QB(n31967) );
  DFFS img_reg_13__1__4_ ( .D(n13160), .CK(clk), .Q(img[372]), .QB(n31954) );
  DFFS img_reg_13__0__4_ ( .D(n13152), .CK(clk), .Q(img[380]), .QB(n31983) );
  DFFS img_reg_14__14__4_ ( .D(n13392), .CK(clk), .Q(img[140]), .QB(n31951) );
  DFFS img_reg_3__14__4_ ( .D(n11984), .CK(clk), .Q(img[1548]), .QB(n31789) );
  DFFS img_reg_1__14__4_ ( .D(n11728), .CK(clk), .Q(img[1804]), .QB(n31773) );
  DFFS img_reg_13__9__4_ ( .D(n13224), .CK(clk), .Q(img[308]), .QB(n31758) );
  DFFS img_reg_10__9__7_ ( .D(n12837), .CK(clk), .Q(img[695]), .QB(n30063) );
  DFFS img_reg_10__9__6_ ( .D(n12838), .CK(clk), .Q(img[694]), .QB(n30451) );
  DFFS img_reg_10__9__5_ ( .D(n12839), .CK(clk), .Q(img[693]), .QB(n30942) );
  DFFS img_reg_10__9__4_ ( .D(n12840), .CK(clk), .Q(img[692]), .QB(n31767) );
  DFFS img_reg_10__9__3_ ( .D(n12841), .CK(clk), .Q(img[691]), .QB(n31429) );
  DFFS img_reg_10__9__2_ ( .D(n12842), .CK(clk), .Q(img[690]), .QB(n30712) );
  DFFS img_reg_10__9__1_ ( .D(n12843), .CK(clk), .Q(img[689]), .QB(n31227) );
  DFFS img_reg_10__9__0_ ( .D(n12844), .CK(clk), .Q(img[688]), .QB(n31725) );
  DFFS img_reg_10__8__7_ ( .D(n12835), .CK(clk), .Q(img[703]), .QB(n30188) );
  DFFS img_reg_10__8__6_ ( .D(n12834), .CK(clk), .Q(img[702]), .QB(n30306) );
  DFFS img_reg_10__8__5_ ( .D(n12833), .CK(clk), .Q(img[701]), .QB(n30919) );
  DFFS img_reg_10__8__3_ ( .D(n12831), .CK(clk), .Q(img[699]), .QB(n31356) );
  DFFS img_reg_10__8__2_ ( .D(n12830), .CK(clk), .Q(img[698]), .QB(n30772) );
  DFFS img_reg_10__8__1_ ( .D(n12829), .CK(clk), .Q(img[697]), .QB(n31242) );
  DFFS img_reg_10__8__0_ ( .D(n12836), .CK(clk), .Q(img[696]), .QB(n31529) );
  DFFS img_reg_10__7__7_ ( .D(n12821), .CK(clk), .Q(img[711]), .QB(n30189) );
  DFFS img_reg_10__7__6_ ( .D(n12822), .CK(clk), .Q(img[710]), .QB(n30307) );
  DFFS img_reg_10__7__5_ ( .D(n12823), .CK(clk), .Q(img[709]), .QB(n30920) );
  DFFS img_reg_10__7__4_ ( .D(n12824), .CK(clk), .Q(img[708]), .QB(n31829) );
  DFFS img_reg_10__7__3_ ( .D(n12825), .CK(clk), .Q(img[707]), .QB(n31357) );
  DFFS img_reg_10__7__2_ ( .D(n12826), .CK(clk), .Q(img[706]), .QB(n30773) );
  DFFS img_reg_10__7__1_ ( .D(n12827), .CK(clk), .Q(img[705]), .QB(n31241) );
  DFFS img_reg_10__7__0_ ( .D(n12828), .CK(clk), .Q(img[704]), .QB(n31530) );
  DFFS img_reg_10__6__7_ ( .D(n12819), .CK(clk), .Q(img[719]), .QB(n30064) );
  DFFS img_reg_10__6__6_ ( .D(n12818), .CK(clk), .Q(img[718]), .QB(n30452) );
  DFFS img_reg_10__6__4_ ( .D(n12816), .CK(clk), .Q(img[716]), .QB(n31768) );
  DFFS img_reg_10__6__3_ ( .D(n12815), .CK(clk), .Q(img[715]), .QB(n31430) );
  DFFS img_reg_10__6__2_ ( .D(n12814), .CK(clk), .Q(img[714]), .QB(n30713) );
  DFFS img_reg_10__6__1_ ( .D(n12813), .CK(clk), .Q(img[713]), .QB(n31228) );
  DFFS img_reg_10__6__0_ ( .D(n12820), .CK(clk), .Q(img[712]), .QB(n31726) );
  DFFS img_reg_10__5__7_ ( .D(n12805), .CK(clk), .Q(img[727]), .QB(n30236) );
  DFFS img_reg_10__5__6_ ( .D(n12806), .CK(clk), .Q(img[726]), .QB(n30511) );
  DFFS img_reg_10__5__5_ ( .D(n12807), .CK(clk), .Q(img[725]), .QB(n30936) );
  DFFS img_reg_10__5__4_ ( .D(n12808), .CK(clk), .Q(img[724]), .QB(n31912) );
  DFFS img_reg_10__5__3_ ( .D(n12809), .CK(clk), .Q(img[723]), .QB(n31330) );
  DFFS img_reg_10__5__2_ ( .D(n12810), .CK(clk), .Q(img[722]), .QB(n30617) );
  DFFS img_reg_10__5__1_ ( .D(n12811), .CK(clk), .Q(img[721]), .QB(n31145) );
  DFFS img_reg_10__5__0_ ( .D(n12812), .CK(clk), .Q(img[720]), .QB(n31711) );
  DFFS img_reg_10__4__7_ ( .D(n12803), .CK(clk), .Q(img[735]), .QB(n30254) );
  DFFS img_reg_10__4__5_ ( .D(n12801), .CK(clk), .Q(img[733]), .QB(n31010) );
  DFFS img_reg_10__4__4_ ( .D(n12800), .CK(clk), .Q(img[732]), .QB(n31972) );
  DFFS img_reg_10__4__3_ ( .D(n12799), .CK(clk), .Q(img[731]), .QB(n31461) );
  DFFS img_reg_10__4__2_ ( .D(n12798), .CK(clk), .Q(img[730]), .QB(n30736) );
  DFFS img_reg_10__4__1_ ( .D(n12797), .CK(clk), .Q(img[729]), .QB(n31098) );
  DFFS img_reg_10__4__0_ ( .D(n12804), .CK(clk), .Q(img[728]), .QB(n31693) );
  DFFS img_reg_10__3__7_ ( .D(n12789), .CK(clk), .Q(img[743]), .QB(n30126) );
  DFFS img_reg_10__3__6_ ( .D(n12790), .CK(clk), .Q(img[742]), .QB(n30432) );
  DFFS img_reg_10__3__5_ ( .D(n12791), .CK(clk), .Q(img[741]), .QB(n30799) );
  DFFS img_reg_10__3__4_ ( .D(n12792), .CK(clk), .Q(img[740]), .QB(n31920) );
  DFFS img_reg_10__3__3_ ( .D(n12793), .CK(clk), .Q(img[739]), .QB(n31496) );
  DFFS img_reg_10__3__2_ ( .D(n12794), .CK(clk), .Q(img[738]), .QB(n30759) );
  DFFS img_reg_10__3__1_ ( .D(n12795), .CK(clk), .Q(img[737]), .QB(n31117) );
  DFFS img_reg_10__3__0_ ( .D(n12796), .CK(clk), .Q(img[736]), .QB(n31741) );
  DFFS img_reg_10__2__6_ ( .D(n12786), .CK(clk), .Q(img[750]), .QB(n30527) );
  DFFS img_reg_10__2__5_ ( .D(n12785), .CK(clk), .Q(img[749]), .QB(n30857) );
  DFFS img_reg_10__2__4_ ( .D(n12784), .CK(clk), .Q(img[748]), .QB(n31893) );
  DFFS img_reg_10__2__3_ ( .D(n12783), .CK(clk), .Q(img[747]), .QB(n31283) );
  DFFS img_reg_10__2__2_ ( .D(n12782), .CK(clk), .Q(img[746]), .QB(n30622) );
  DFFS img_reg_10__2__1_ ( .D(n12781), .CK(clk), .Q(img[745]), .QB(n31256) );
  DFFS img_reg_10__2__0_ ( .D(n12788), .CK(clk), .Q(img[744]), .QB(n31599) );
  DFFS img_reg_10__1__7_ ( .D(n12773), .CK(clk), .Q(img[759]), .QB(n30267) );
  DFFS img_reg_10__1__6_ ( .D(n12774), .CK(clk), .Q(img[758]), .QB(n30370) );
  DFFS img_reg_10__1__5_ ( .D(n12775), .CK(clk), .Q(img[757]), .QB(n30981) );
  DFFS img_reg_10__1__4_ ( .D(n12776), .CK(clk), .Q(img[756]), .QB(n31959) );
  DFFS img_reg_10__1__3_ ( .D(n12777), .CK(clk), .Q(img[755]), .QB(n31413) );
  DFFS img_reg_10__1__2_ ( .D(n12778), .CK(clk), .Q(img[754]), .QB(n30553) );
  DFFS img_reg_10__1__1_ ( .D(n12779), .CK(clk), .Q(img[753]), .QB(n31206) );
  DFFS img_reg_10__0__7_ ( .D(n12771), .CK(clk), .Q(img[767]), .QB(n30281) );
  DFFS img_reg_10__0__6_ ( .D(n12770), .CK(clk), .Q(img[766]), .QB(n30481) );
  DFFS img_reg_10__0__5_ ( .D(n12769), .CK(clk), .Q(img[765]), .QB(n30995) );
  DFFS img_reg_10__0__4_ ( .D(n12768), .CK(clk), .Q(img[764]), .QB(n31987) );
  DFFS img_reg_10__0__3_ ( .D(n12767), .CK(clk), .Q(img[763]), .QB(n31480) );
  DFFS img_reg_10__0__2_ ( .D(n12766), .CK(clk), .Q(img[762]), .QB(n30666) );
  DFFS img_reg_10__0__1_ ( .D(n12765), .CK(clk), .Q(img[761]), .QB(n31036) );
  DFFS img_reg_10__0__0_ ( .D(n12772), .CK(clk), .Q(img[760]), .QB(n31571) );
  DFFS img_reg_0__11__7_ ( .D(n11573), .CK(clk), .Q(img[1959]), .QB(n30160) );
  DFFS img_reg_0__11__6_ ( .D(n11574), .CK(clk), .Q(img[1958]), .QB(n30336) );
  DFFS img_reg_0__11__5_ ( .D(n11575), .CK(clk), .Q(img[1957]), .QB(n30828) );
  DFFS img_reg_0__11__4_ ( .D(n11576), .CK(clk), .Q(img[1956]), .QB(n31859) );
  DFFS img_reg_0__11__3_ ( .D(n11577), .CK(clk), .Q(img[1955]), .QB(n31383) );
  DFFS img_reg_0__11__2_ ( .D(n11578), .CK(clk), .Q(img[1954]), .QB(n30641) );
  DFFS img_reg_0__11__0_ ( .D(n11580), .CK(clk), .Q(img[1952]), .QB(n31551) );
  DFFS img_reg_2__11__7_ ( .D(n11829), .CK(clk), .Q(img[1703]), .QB(n30140) );
  DFFS img_reg_2__11__6_ ( .D(n11830), .CK(clk), .Q(img[1702]), .QB(n30316) );
  DFFS img_reg_2__11__5_ ( .D(n11831), .CK(clk), .Q(img[1701]), .QB(n30810) );
  DFFS img_reg_2__11__4_ ( .D(n11832), .CK(clk), .Q(img[1700]), .QB(n31839) );
  DFFS img_reg_2__11__3_ ( .D(n11833), .CK(clk), .Q(img[1699]), .QB(n31366) );
  DFFS img_reg_2__11__2_ ( .D(n11834), .CK(clk), .Q(img[1698]), .QB(n30675) );
  DFFS img_reg_2__11__1_ ( .D(n11835), .CK(clk), .Q(img[1697]), .QB(n31046) );
  DFFS img_reg_2__11__0_ ( .D(n11836), .CK(clk), .Q(img[1696]), .QB(n31531) );
  DFFS img_reg_11__11__7_ ( .D(n12985), .CK(clk), .Q(img[551]), .QB(n30242) );
  DFFS img_reg_11__11__6_ ( .D(n12984), .CK(clk), .Q(img[550]), .QB(n30453) );
  DFFS img_reg_11__11__5_ ( .D(n12983), .CK(clk), .Q(img[549]), .QB(n31992) );
  DFFS img_reg_11__11__4_ ( .D(n12982), .CK(clk), .Q(img[548]), .QB(n31960) );
  DFFS img_reg_11__11__3_ ( .D(n12981), .CK(clk), .Q(img[547]), .QB(n31990) );
  DFFS img_reg_11__11__1_ ( .D(n12987), .CK(clk), .Q(img[545]), .QB(n31074) );
  DFFS img_reg_11__11__0_ ( .D(n12988), .CK(clk), .Q(img[544]), .QB(n31667) );
  DFFS img_reg_2__4__2_ ( .D(n11774), .CK(clk), .Q(img[1754]), .QB(n30676) );
  DFFS img_reg_1__4__2_ ( .D(n11650), .CK(clk), .Q(img[1882]), .QB(n30668) );
  DFFS img_reg_1__4__0_ ( .D(n11652), .CK(clk), .Q(img[1880]), .QB(n31502) );
  QDFFS img_reg_9__6__4_ ( .D(n12688), .CK(clk), .Q(img[844]) );
  QDFFS img_reg_0__6__5_ ( .D(n11537), .CK(clk), .Q(img[1997]) );
  DFFS img_reg_0__7__7_ ( .D(n11541), .CK(clk), .Q(img[1991]), .QB(n30157) );
  DFFS img_reg_5__3__6_ ( .D(n12154), .CK(clk), .Q(img[1382]), .QB(n30417) );
  DFFS img_reg_2__0__1_ ( .D(n11741), .CK(clk), .Q(img[1785]), .QB(n31052) );
  DFFS img_reg_5__0__4_ ( .D(n12128), .CK(clk), .Q(img[1404]), .QB(n31814) );
  DFFS img_reg_4__5__5_ ( .D(n12039), .CK(clk), .Q(img[1493]), .QB(n30853) );
  DFFS img_reg_5__6__5_ ( .D(n12175), .CK(clk), .Q(img[1357]), .QB(n30954) );
  DFFS img_reg_2__1__5_ ( .D(n11751), .CK(clk), .Q(img[1781]), .QB(n30870) );
  DFFS img_reg_3__0__5_ ( .D(n11871), .CK(clk), .Q(img[1661]), .QB(n30816) );
  DFFS img_reg_7__5__0_ ( .D(n12428), .CK(clk), .Q(img[1104]), .QB(n31625) );
  DFFS img_reg_2__7__0_ ( .D(n11804), .CK(clk), .Q(img[1728]), .QB(n31538) );
  DFFS img_reg_5__0__0_ ( .D(n12132), .CK(clk), .Q(img[1400]), .QB(n31518) );
  DFFS img_reg_6__3__0_ ( .D(n12284), .CK(clk), .Q(img[1248]), .QB(n31672) );
  DFFS img_reg_3__0__2_ ( .D(n11874), .CK(clk), .Q(img[1658]), .QB(n30690) );
  DFFS img_reg_5__5__3_ ( .D(n12167), .CK(clk), .Q(img[1363]), .QB(n31267) );
  DFFS img_reg_5__1__3_ ( .D(n12135), .CK(clk), .Q(img[1395]), .QB(n31399) );
  DFFS img_reg_1__0__3_ ( .D(n11617), .CK(clk), .Q(img[1915]), .QB(n31363) );
  DFFS img_reg_6__5__1_ ( .D(n12299), .CK(clk), .Q(img[1233]), .QB(n31126) );
  DFFS img_reg_7__3__1_ ( .D(n12405), .CK(clk), .Q(img[1121]), .QB(n31101) );
  DFFS img_reg_5__2__6_ ( .D(n12142), .CK(clk), .Q(img[1390]), .QB(n30483) );
  DFFS img_reg_6__2__6_ ( .D(n12274), .CK(clk), .Q(img[1262]), .QB(n30499) );
  DFFS img_reg_2__6__7_ ( .D(n11795), .CK(clk), .Q(img[1743]), .QB(n30080) );
  DFFS img_reg_5__2__7_ ( .D(n12141), .CK(clk), .Q(img[1391]), .QB(n30204) );
  DFFS img_reg_1__0__1_ ( .D(n11619), .CK(clk), .Q(img[1913]), .QB(n31044) );
  DFFS img_reg_0__3__6_ ( .D(n11510), .CK(clk), .Q(img[2022]), .QB(n30339) );
  DFFS img_reg_2__6__4_ ( .D(n11792), .CK(clk), .Q(img[1740]), .QB(n31784) );
  DFFS img_reg_6__3__4_ ( .D(n12280), .CK(clk), .Q(img[1252]), .QB(n31924) );
  DFFS img_reg_2__2__4_ ( .D(n11760), .CK(clk), .Q(img[1772]), .QB(n31780) );
  DFFS img_reg_15__8__5_ ( .D(n13471), .CK(clk), .Q(img[61]), .QB(n30896) );
  DFFS img_reg_3__13__0_ ( .D(n11980), .CK(clk), .Q(img[1552]), .QB(n31622) );
  DFFS img_reg_14__15__5_ ( .D(n13399), .CK(clk), .Q(img[133]), .QB(n30982) );
  DFFS img_reg_5__12__5_ ( .D(n12223), .CK(clk), .Q(img[1309]), .QB(n30784) );
  DFFS img_reg_1__8__5_ ( .D(n11679), .CK(clk), .Q(img[1853]), .QB(n30800) );
  DFFS img_reg_9__12__5_ ( .D(n12735), .CK(clk), .Q(img[797]), .QB(n30797) );
  DFFS img_reg_11__5__5_ ( .D(n12937), .CK(clk), .Q(img[597]), .QB(n30922) );
  DFFS img_reg_11__9__2_ ( .D(n12966), .CK(clk), .Q(img[562]), .QB(n30699) );
  DFFS img_reg_5__11__3_ ( .D(n12215), .CK(clk), .Q(img[1315]), .QB(n31450) );
  DFFS img_reg_5__13__3_ ( .D(n12231), .CK(clk), .Q(img[1299]), .QB(n31269) );
  DFFS img_reg_14__2__3_ ( .D(n13295), .CK(clk), .Q(img[235]), .QB(n31272) );
  DFFS img_reg_12__5__3_ ( .D(n13065), .CK(clk), .Q(img[467]), .QB(n31326) );
  DFFS img_reg_6__8__3_ ( .D(n12319), .CK(clk), .Q(img[1211]), .QB(n31338) );
  DFFS img_reg_8__2__4_ ( .D(n12528), .CK(clk), .Q(img[1004]), .QB(n31880) );
  DFFS img_reg_11__7__2_ ( .D(n12950), .CK(clk), .Q(img[578]), .QB(n30761) );
  DFFS img_reg_5__13__0_ ( .D(n12236), .CK(clk), .Q(img[1296]), .QB(n31583) );
  DFFS img_reg_14__2__0_ ( .D(n13300), .CK(clk), .Q(img[232]), .QB(n31588) );
  DFFS img_reg_14__6__2_ ( .D(n13326), .CK(clk), .Q(img[202]), .QB(n30706) );
  DFFS img_reg_14__0__0_ ( .D(n13284), .CK(clk), .Q(img[248]), .QB(n31565) );
  DFFS img_reg_6__8__2_ ( .D(n12318), .CK(clk), .Q(img[1210]), .QB(n30637) );
  DFFS img_reg_11__8__1_ ( .D(n12963), .CK(clk), .Q(img[569]), .QB(n31230) );
  DFFS img_reg_5__13__1_ ( .D(n12229), .CK(clk), .Q(img[1297]), .QB(n31127) );
  DFFS img_reg_14__9__6_ ( .D(n13350), .CK(clk), .Q(img[182]), .QB(n30444) );
  DFFS img_reg_14__6__1_ ( .D(n13325), .CK(clk), .Q(img[201]), .QB(n31220) );
  DFFS img_reg_12__2__6_ ( .D(n13042), .CK(clk), .Q(img[494]), .QB(n30524) );
  DFFS img_reg_3__10__7_ ( .D(n11949), .CK(clk), .Q(img[1583]), .QB(n30081) );
  DFFS img_reg_5__13__7_ ( .D(n12235), .CK(clk), .Q(img[1303]), .QB(n30205) );
  DFFS img_reg_14__10__7_ ( .D(n13363), .CK(clk), .Q(img[175]), .QB(n30230) );
  DFFS img_reg_0__8__7_ ( .D(n11555), .CK(clk), .Q(img[1983]), .QB(n30156) );
  DFFS img_reg_4__12__4_ ( .D(n12096), .CK(clk), .Q(img[1436]), .QB(n31935) );
  DFFS img_reg_0__13__4_ ( .D(n11592), .CK(clk), .Q(img[1940]), .QB(n31799) );
  DFFS img_reg_0__12__4_ ( .D(n11584), .CK(clk), .Q(img[1948]), .QB(n31861) );
  DFFS img_reg_12__4__4_ ( .D(n13056), .CK(clk), .Q(img[476]), .QB(n31969) );
  DFFS img_reg_15__0__4_ ( .D(n13408), .CK(clk), .Q(img[124]), .QB(n31977) );
  DFFS img_reg_5__6__0_ ( .D(n12180), .CK(clk), .Q(img[1352]), .QB(n31645) );
  DFFS img_reg_1__7__2_ ( .D(n11670), .CK(clk), .Q(img[1858]), .QB(n30672) );
  QDFFN img_reg_5__0__5_ ( .D(n12127), .CK(clk), .Q(img[1405]) );
  QDFFN img_reg_9__5__4_ ( .D(n12680), .CK(clk), .Q(img[852]) );
  QDFFN img_reg_9__2__4_ ( .D(n12656), .CK(clk), .Q(img[876]) );
  QDFFN img_reg_9__3__5_ ( .D(n12665), .CK(clk), .Q(img[869]) );
  QDFFN img_reg_9__2__5_ ( .D(n12655), .CK(clk), .Q(img[877]) );
  QDFFN img_reg_9__7__5_ ( .D(n12697), .CK(clk), .Q(img[837]) );
  QDFFN img_reg_9__1__4_ ( .D(n12648), .CK(clk), .Q(img[884]) );
  QDFFN img_reg_9__0__5_ ( .D(n12639), .CK(clk), .Q(img[893]) );
  QDFFN img_reg_12__0__4_ ( .D(n13024), .CK(clk), .Q(img[508]) );
  QDFFN img_reg_1__4__5_ ( .D(n11647), .CK(clk), .Q(img[1885]) );
  QDFFN img_reg_9__0__4_ ( .D(n12640), .CK(clk), .Q(img[892]) );
  QDFFN img_reg_12__0__5_ ( .D(n13025), .CK(clk), .Q(img[509]) );
  QDFFN img_reg_9__7__4_ ( .D(n12696), .CK(clk), .Q(img[836]) );
  QDFFN img_reg_1__7__5_ ( .D(n11673), .CK(clk), .Q(img[1861]) );
  QDFFN img_reg_6__0__5_ ( .D(n12257), .CK(clk), .Q(img[1277]) );
  QDFFN img_reg_6__7__5_ ( .D(n12311), .CK(clk), .Q(img[1221]) );
  OAI12HS U13755 ( .B1(n24023), .B2(n24466), .A1(n24495), .O(n29040) );
  INV1S U13756 ( .I(n23380), .O(n23387) );
  OAI12HS U13757 ( .B1(n22860), .B2(n22810), .A1(n22809), .O(n22855) );
  AOI13HS U13758 ( .B1(n29518), .B2(n29469), .B3(n29516), .A1(n29468), .O(
        n29473) );
  AOI12HS U13759 ( .B1(n22768), .B2(n22872), .A1(n22767), .O(n22860) );
  INV1S U13760 ( .I(n24203), .O(n24669) );
  MOAI1S U13761 ( .A1(n28573), .A2(n27914), .B1(n28571), .B2(n27913), .O(
        n27915) );
  NR2P U13762 ( .I1(n23915), .I2(n24098), .O(n24463) );
  OAI12HS U13763 ( .B1(n28536), .B2(n27266), .A1(n27265), .O(n27289) );
  OAI12HS U13764 ( .B1(n28536), .B2(n25395), .A1(n25394), .O(n25420) );
  OAI12HS U13765 ( .B1(n28536), .B2(n21624), .A1(n28535), .O(n28576) );
  NR2 U13766 ( .I1(n24002), .I2(n24013), .O(n24673) );
  NR2 U13767 ( .I1(n23284), .I2(n23285), .O(n23389) );
  AOI12HS U13768 ( .B1(n28534), .B2(n28533), .A1(n28532), .O(n28535) );
  AOI12HS U13769 ( .B1(n28534), .B2(n29443), .A1(n27264), .O(n27265) );
  OR2 U13770 ( .I1(n24706), .I2(n13908), .O(n28573) );
  AOI12HS U13771 ( .B1(n28534), .B2(n29505), .A1(n24770), .O(n24771) );
  BUF1 U13772 ( .I(n21456), .O(n29507) );
  OA12 U13773 ( .B1(n24699), .B2(n23898), .A1(n23956), .O(n24722) );
  FA1S U13774 ( .A(n22375), .B(n22374), .CI(n22373), .CO(n22403), .S(n22377)
         );
  FA1S U13775 ( .A(n22372), .B(n22371), .CI(n22370), .CO(n22392), .S(n22394)
         );
  OR2 U13776 ( .I1(n23893), .I2(n23894), .O(n24700) );
  INV1S U13777 ( .I(n20668), .O(n20669) );
  FA1S U13778 ( .A(n21668), .B(n21667), .CI(n21666), .CO(n22369), .S(n21685)
         );
  FA1S U13779 ( .A(n21682), .B(n21681), .CI(n21680), .CO(n21664), .S(n21699)
         );
  FA1S U13780 ( .A(n21698), .B(n21697), .CI(n21696), .CO(n21720), .S(n22383)
         );
  OR2 U13781 ( .I1(n23895), .I2(n23894), .O(n24699) );
  INV2 U13782 ( .I(n22410), .O(n22523) );
  FA1S U13783 ( .A(n21775), .B(n21774), .CI(n21773), .CO(n21801), .S(n21777)
         );
  NR2 U13784 ( .I1(n29968), .I2(n13822), .O(n23770) );
  INV1S U13785 ( .I(n21374), .O(n21379) );
  INV1S U13786 ( .I(n30029), .O(n23640) );
  FA1S U13787 ( .A(n22390), .B(n22389), .CI(n22388), .CO(n22386), .S(PE_N82)
         );
  FA1S U13788 ( .A(n21695), .B(n21694), .CI(n21693), .CO(n21696), .S(n22385)
         );
  INV1S U13789 ( .I(n23179), .O(n23297) );
  FA1S U13790 ( .A(n21769), .B(n21768), .CI(n21767), .CO(n21797), .S(n21773)
         );
  FA1S U13791 ( .A(n15926), .B(n15925), .CI(n15924), .CO(n15941), .S(n15952)
         );
  OAI12HP U13792 ( .B1(n21104), .B2(n21103), .A1(n21109), .O(n23841) );
  AO12P U13793 ( .B1(n19441), .B2(n19440), .A1(n19439), .O(n21472) );
  ND2P U13794 ( .I1(n21092), .I2(n21091), .O(n21109) );
  INV1S U13795 ( .I(n20921), .O(n20840) );
  OA112 U13796 ( .C1(n13818), .C2(n22941), .A1(n22935), .B1(n22934), .O(n22936) );
  INV1S U13797 ( .I(n30027), .O(n23559) );
  FA1S U13798 ( .A(n15894), .B(n15893), .CI(n15892), .CO(n15895), .S(n21764)
         );
  AO12 U13799 ( .B1(n20791), .B2(n20790), .A1(n20789), .O(n13909) );
  INV1S U13800 ( .I(n21194), .O(n21206) );
  INV1S U13801 ( .I(n21812), .O(n21849) );
  FA1S U13802 ( .A(n15855), .B(n15854), .CI(n15853), .CO(n21784), .S(n21785)
         );
  FA1S U13803 ( .A(n21790), .B(n21789), .CI(n21788), .CO(n21786), .S(PE_N50)
         );
  INV1S U13804 ( .I(n20605), .O(n21729) );
  INV2 U13805 ( .I(n21088), .O(n29505) );
  INV3 U13806 ( .I(n22059), .O(n22162) );
  ND2 U13807 ( .I1(n21669), .I2(n20809), .O(n20788) );
  AOI12HS U13808 ( .B1(n16260), .B2(n19533), .A1(n16259), .O(n16261) );
  ND3 U13809 ( .I1(n16214), .I2(n16213), .I3(n16215), .O(n21803) );
  ND2 U13810 ( .I1(n21653), .I2(n20809), .O(n20784) );
  NR2T U13811 ( .I1(n21345), .I2(n20601), .O(n29509) );
  INV2 U13812 ( .I(n20863), .O(n13817) );
  AO12P U13813 ( .B1(n20568), .B2(n20567), .A1(n21340), .O(n26013) );
  INV1S U13814 ( .I(n21616), .O(n21656) );
  ND3P U13815 ( .I1(n20290), .I2(n20289), .I3(n20288), .O(n22661) );
  NR2P U13816 ( .I1(n13822), .I2(n20605), .O(n21345) );
  NR2P U13817 ( .I1(n13822), .I2(n20537), .O(n21340) );
  BUF3 U13818 ( .I(n21398), .O(n29497) );
  ND3P U13819 ( .I1(n17435), .I2(n17434), .I3(n17433), .O(n22058) );
  NR2 U13820 ( .I1(n13822), .I2(n21236), .O(n21346) );
  INV2 U13821 ( .I(n22932), .O(n13816) );
  NR2P U13822 ( .I1(n13822), .I2(n20436), .O(n21330) );
  OR2 U13823 ( .I1(n13822), .I2(n23180), .O(n21000) );
  ND2 U13824 ( .I1(n19227), .I2(n19226), .O(n19232) );
  OR2P U13825 ( .I1(n19706), .I2(n19705), .O(n23185) );
  ND2 U13826 ( .I1(n16026), .I2(n16025), .O(n20610) );
  ND2 U13827 ( .I1(n16015), .I2(n16014), .O(n20611) );
  ND2 U13828 ( .I1(n16199), .I2(n16198), .O(n20608) );
  MXL2H U13829 ( .A(n22667), .B(n20358), .S(n13822), .OB(n25391) );
  ND2 U13830 ( .I1(n16273), .I2(n16272), .O(n20593) );
  ND2 U13831 ( .I1(n16381), .I2(n16380), .O(n20585) );
  ND2 U13832 ( .I1(n16359), .I2(n16358), .O(n20595) );
  ND2 U13833 ( .I1(n19277), .I2(n19276), .O(n20233) );
  ND2 U13834 ( .I1(n16336), .I2(n16335), .O(n20573) );
  ND2 U13835 ( .I1(n16325), .I2(n16324), .O(n20570) );
  ND2 U13836 ( .I1(n16651), .I2(n16650), .O(n20561) );
  ND2 U13837 ( .I1(n16566), .I2(n16565), .O(n20552) );
  ND2 U13838 ( .I1(n16536), .I2(n16535), .O(n20551) );
  ND2S U13839 ( .I1(n19513), .I2(n19512), .O(n19519) );
  ND2 U13840 ( .I1(n19968), .I2(n19967), .O(n20298) );
  ND2 U13841 ( .I1(n16620), .I2(n16619), .O(n20539) );
  ND2 U13842 ( .I1(n16514), .I2(n16513), .O(n20544) );
  ND2 U13843 ( .I1(n16401), .I2(n16400), .O(n19929) );
  ND2 U13844 ( .I1(n16600), .I2(n16599), .O(n20546) );
  ND2 U13845 ( .I1(n16641), .I2(n16640), .O(n20013) );
  ND2 U13846 ( .I1(n16610), .I2(n16609), .O(n20558) );
  ND2 U13847 ( .I1(n17740), .I2(n17739), .O(n20511) );
  ND2 U13848 ( .I1(n17718), .I2(n17717), .O(n20513) );
  ND2 U13849 ( .I1(n17761), .I2(n17760), .O(n20507) );
  AOI12HS U13850 ( .B1(n20350), .B2(n20364), .A1(n20349), .O(n20353) );
  ND2 U13851 ( .I1(n17856), .I2(n17855), .O(n20522) );
  ND2 U13852 ( .I1(n17846), .I2(n17845), .O(n20527) );
  ND2 U13853 ( .I1(n17728), .I2(n17727), .O(n20526) );
  ND2 U13854 ( .I1(n17707), .I2(n17706), .O(n20512) );
  ND2 U13855 ( .I1(n17834), .I2(n17833), .O(n20520) );
  AOI22S U13856 ( .A1(n20350), .A2(n20371), .B1(n20363), .B2(n20350), .O(
        n20354) );
  ND2 U13857 ( .I1(n18952), .I2(n18951), .O(n20075) );
  ND2 U13858 ( .I1(n17822), .I2(n17821), .O(n20508) );
  ND2 U13859 ( .I1(n17809), .I2(n17808), .O(n20521) );
  ND2 U13860 ( .I1(n18929), .I2(n18928), .O(n20084) );
  ND2 U13861 ( .I1(n18879), .I2(n18878), .O(n20069) );
  ND2 U13862 ( .I1(n17799), .I2(n17798), .O(n20514) );
  ND2 U13863 ( .I1(n19030), .I2(n19029), .O(n20086) );
  ND2 U13864 ( .I1(n18969), .I2(n18968), .O(n20073) );
  ND2 U13865 ( .I1(n18891), .I2(n18890), .O(n20072) );
  ND2 U13866 ( .I1(n17270), .I2(n17269), .O(n20490) );
  ND2 U13867 ( .I1(n18104), .I2(n18103), .O(n20334) );
  ND2 U13868 ( .I1(n17567), .I2(n17566), .O(n20428) );
  ND2 U13869 ( .I1(n17577), .I2(n17576), .O(n20403) );
  OAI112HS U13870 ( .C1(n16713), .C2(n15142), .A1(n15036), .B1(n15035), .O(
        n15037) );
  OR2P U13871 ( .I1(n18133), .I2(n19700), .O(n19542) );
  NR2 U13872 ( .I1(n20969), .I2(n14503), .O(n19534) );
  ND2 U13873 ( .I1(n16764), .I2(n16763), .O(n20445) );
  ND2 U13874 ( .I1(n16805), .I2(n16804), .O(n20437) );
  ND2 U13875 ( .I1(n16774), .I2(n16773), .O(n20457) );
  ND2 U13876 ( .I1(n16815), .I2(n16814), .O(n20456) );
  ND2S U13877 ( .I1(n19092), .I2(n19091), .O(n19983) );
  ND2 U13878 ( .I1(n16825), .I2(n16824), .O(n20455) );
  ND2 U13879 ( .I1(n16869), .I2(n16868), .O(n20452) );
  AN4S U13880 ( .I1(n17597), .I2(n17596), .I3(n17595), .I4(n17594), .O(n17598)
         );
  AN4S U13881 ( .I1(n17608), .I2(n17607), .I3(n17606), .I4(n17605), .O(n17609)
         );
  ND2 U13882 ( .I1(n17125), .I2(n17124), .O(n21038) );
  ND2 U13883 ( .I1(n17207), .I2(n17206), .O(n20471) );
  ND2 U13884 ( .I1(n16879), .I2(n16878), .O(n20458) );
  ND2 U13885 ( .I1(n17009), .I2(n17008), .O(n21040) );
  ND2 U13886 ( .I1(n17228), .I2(n17227), .O(n20492) );
  ND2 U13887 ( .I1(n17114), .I2(n17113), .O(n21063) );
  ND2 U13888 ( .I1(n16989), .I2(n16988), .O(n21043) );
  ND2 U13889 ( .I1(n17029), .I2(n17028), .O(n21050) );
  ND2 U13890 ( .I1(n16999), .I2(n16998), .O(n21049) );
  ND2 U13891 ( .I1(n17019), .I2(n17018), .O(n21058) );
  ND2 U13892 ( .I1(n16794), .I2(n16793), .O(n20451) );
  ND2 U13893 ( .I1(n16784), .I2(n16783), .O(n20443) );
  ND2 U13894 ( .I1(n17297), .I2(n17296), .O(n20468) );
  ND2 U13895 ( .I1(n17083), .I2(n17082), .O(n21037) );
  ND2 U13896 ( .I1(n17094), .I2(n17093), .O(n21046) );
  ND2 U13897 ( .I1(n16859), .I2(n16858), .O(n20440) );
  ND2 U13898 ( .I1(n18457), .I2(n18456), .O(n20344) );
  ND2 U13899 ( .I1(n19199), .I2(n19198), .O(n20293) );
  ND2 U13900 ( .I1(n17353), .I2(n17352), .O(n20476) );
  ND2 U13901 ( .I1(n17329), .I2(n17328), .O(n20475) );
  ND2 U13902 ( .I1(n17217), .I2(n17216), .O(n20489) );
  ND2 U13903 ( .I1(n17260), .I2(n17259), .O(n20485) );
  ND2 U13904 ( .I1(n16753), .I2(n16752), .O(n20444) );
  ND2 U13905 ( .I1(n17533), .I2(n17532), .O(n20419) );
  ND2 U13906 ( .I1(n17521), .I2(n17520), .O(n20404) );
  MOAI1S U13907 ( .A1(n17414), .A2(n13929), .B1(n17413), .B2(n13839), .O(
        n14436) );
  AN4S U13908 ( .I1(n16823), .I2(n16822), .I3(n16821), .I4(n16820), .O(n16824)
         );
  AN4S U13909 ( .I1(n17061), .I2(n17060), .I3(n17059), .I4(n17058), .O(n17062)
         );
  AN4S U13910 ( .I1(n16887), .I2(n16886), .I3(n16885), .I4(n16884), .O(n16888)
         );
  MOAI1S U13911 ( .A1(n16935), .A2(n17656), .B1(n16934), .B2(n17931), .O(
        n16936) );
  AN4S U13912 ( .I1(n16837), .I2(n16836), .I3(n16835), .I4(n16834), .O(n16838)
         );
  ND2S U13913 ( .I1(n18784), .I2(n18783), .O(n20143) );
  ND2S U13914 ( .I1(n18771), .I2(n18770), .O(n20153) );
  ND2 U13915 ( .I1(n18349), .I2(n18348), .O(n19835) );
  ND2 U13916 ( .I1(n18523), .I2(n18522), .O(n19754) );
  ND2 U13917 ( .I1(n18691), .I2(n18690), .O(n20139) );
  ND2S U13918 ( .I1(n18381), .I2(n18380), .O(n19827) );
  ND2S U13919 ( .I1(n18598), .I2(n18597), .O(n19755) );
  ND2S U13920 ( .I1(n18807), .I2(n18806), .O(n20141) );
  ND2S U13921 ( .I1(n18830), .I2(n18829), .O(n20154) );
  ND2 U13922 ( .I1(n18608), .I2(n18607), .O(n19743) );
  ND2S U13923 ( .I1(n18533), .I2(n18532), .O(n19758) );
  ND2S U13924 ( .I1(n18712), .I2(n18711), .O(n20142) );
  ND2S U13925 ( .I1(n18757), .I2(n18756), .O(n20140) );
  ND2S U13926 ( .I1(n18795), .I2(n18794), .O(n20152) );
  ND2 U13927 ( .I1(n18503), .I2(n18502), .O(n19770) );
  ND2 U13928 ( .I1(n18680), .I2(n18679), .O(n20163) );
  ND2 U13929 ( .I1(n18574), .I2(n18573), .O(n19752) );
  ND2 U13930 ( .I1(n18175), .I2(n18174), .O(n19684) );
  AN4S U13931 ( .I1(n17102), .I2(n17101), .I3(n17100), .I4(n17099), .O(n17103)
         );
  ND2 U13932 ( .I1(n18185), .I2(n18184), .O(n19674) );
  ND2 U13933 ( .I1(n18329), .I2(n18328), .O(n19837) );
  ND2 U13934 ( .I1(n18639), .I2(n18638), .O(n19742) );
  ND2 U13935 ( .I1(n18543), .I2(n18542), .O(n19756) );
  NR2 U13936 ( .I1(n15302), .I2(n15301), .O(n15354) );
  NR2 U13937 ( .I1(n15772), .I2(n15771), .O(n16233) );
  AN4S U13938 ( .I1(n18205), .I2(n18204), .I3(n18203), .I4(n18202), .O(n18206)
         );
  AN4S U13939 ( .I1(n18782), .I2(n18781), .I3(n18780), .I4(n18779), .O(n18783)
         );
  AN4S U13940 ( .I1(n18765), .I2(n18764), .I3(n18763), .I4(n18762), .O(n18771)
         );
  AN4S U13941 ( .I1(n18815), .I2(n18814), .I3(n18813), .I4(n18812), .O(n18816)
         );
  AN4S U13942 ( .I1(n18572), .I2(n18571), .I3(n18570), .I4(n18569), .O(n18573)
         );
  NR2 U13943 ( .I1(n14952), .I2(n14951), .O(n16706) );
  NR2 U13944 ( .I1(n14978), .I2(n14977), .O(n16708) );
  NR2 U13945 ( .I1(n15001), .I2(n15000), .O(n16713) );
  AN4S U13946 ( .I1(n18183), .I2(n18182), .I3(n18181), .I4(n18180), .O(n18184)
         );
  NR2 U13947 ( .I1(n15511), .I2(n15510), .O(n16482) );
  ND3 U13948 ( .I1(n15522), .I2(n15521), .I3(n15520), .O(n16476) );
  NR2 U13949 ( .I1(n15390), .I2(n15389), .O(n16471) );
  AOI22S U13950 ( .A1(n17404), .A2(n13847), .B1(n21062), .B2(n17403), .O(
        n14383) );
  MOAI1S U13951 ( .A1(n16946), .A2(n15142), .B1(n16945), .B2(n18040), .O(
        n14282) );
  AN4S U13952 ( .I1(n15394), .I2(n15393), .I3(n15392), .I4(n15391), .O(n15401)
         );
  AN4S U13953 ( .I1(n14982), .I2(n14981), .I3(n14980), .I4(n14979), .O(n14989)
         );
  AN4S U13954 ( .I1(n15079), .I2(n15078), .I3(n15077), .I4(n15076), .O(n15087)
         );
  NR2 U13955 ( .I1(n14399), .I2(n14398), .O(n17412) );
  NR2 U13956 ( .I1(n14733), .I2(n14732), .O(n17657) );
  NR2 U13957 ( .I1(n14472), .I2(n14471), .O(n17421) );
  NR2 U13958 ( .I1(n14758), .I2(n14757), .O(n17659) );
  NR2 U13959 ( .I1(n15265), .I2(n15264), .O(n17930) );
  INV2 U13960 ( .I(n20421), .O(n18040) );
  BUF2 U13961 ( .I(n14739), .O(n13798) );
  AN4S U13962 ( .I1(n14861), .I2(n14860), .I3(n14859), .I4(n14858), .O(n14868)
         );
  NR2 U13963 ( .I1(n14666), .I2(n14665), .O(n17164) );
  NR2 U13964 ( .I1(n14689), .I2(n14688), .O(n17159) );
  NR2 U13965 ( .I1(n14424), .I2(n14423), .O(n17414) );
  NR2 U13966 ( .I1(n14186), .I2(n14185), .O(n16933) );
  NR2 U13967 ( .I1(n14089), .I2(n14088), .O(n16946) );
  NR2 U13968 ( .I1(n14449), .I2(n14448), .O(n17417) );
  NR2 U13969 ( .I1(n14172), .I2(n14171), .O(n16954) );
  ND2 U13970 ( .I1(n23835), .I2(n14105), .O(n20421) );
  BUF4 U13971 ( .I(n14822), .O(n18946) );
  BUF2 U13972 ( .I(n16353), .O(n17827) );
  BUF2 U13973 ( .I(n13803), .O(n17778) );
  BUF2 U13974 ( .I(n18148), .O(n18911) );
  BUF2 U13975 ( .I(n13803), .O(n18996) );
  BUF3 U13976 ( .I(n15568), .O(n19326) );
  INV3 U13977 ( .I(n17522), .O(n16048) );
  BUF6 U13978 ( .I(n13827), .O(n13783) );
  INV2 U13979 ( .I(n28540), .O(n28555) );
  INV3 U13980 ( .I(n18297), .O(n19023) );
  NR2P U13981 ( .I1(n23642), .I2(act_ptr[1]), .O(n13989) );
  BUF1 U13982 ( .I(n19245), .O(n18837) );
  NR2P U13983 ( .I1(n23642), .I2(n13959), .O(n13986) );
  BUF2 U13984 ( .I(n13886), .O(n13875) );
  BUF2 U13985 ( .I(n14822), .O(n16515) );
  NR2P U13986 ( .I1(n23900), .I2(n23973), .O(n23954) );
  BUF4 U13987 ( .I(n17515), .O(n13841) );
  BUF8CK U13988 ( .I(n13931), .O(n13845) );
  INV6 U13989 ( .I(n15277), .O(n15568) );
  BUF4 U13990 ( .I(n15752), .O(n13885) );
  BUF4 U13991 ( .I(n15752), .O(n13884) );
  INV1S U13992 ( .I(n19024), .O(n13873) );
  INV2 U13993 ( .I(n20191), .O(n13857) );
  BUF4 U13994 ( .I(n18155), .O(n13886) );
  BUF1 U13995 ( .I(n13840), .O(n15801) );
  BUF2 U13996 ( .I(n13931), .O(n14739) );
  BUF3 U13997 ( .I(n16002), .O(n13848) );
  BUF6CK U13998 ( .I(n16003), .O(n17880) );
  INV6 U13999 ( .I(n17886), .O(n15674) );
  INV2 U14000 ( .I(n16326), .O(n13834) );
  INV3CK U14001 ( .I(n16003), .O(n14034) );
  INV1 U14002 ( .I(n14077), .O(n16431) );
  NR2P U14003 ( .I1(i_row[0]), .I2(n14043), .O(n14045) );
  BUF2 U14004 ( .I(n16375), .O(n14299) );
  ND2T U14005 ( .I1(i_row[1]), .I2(i_row[2]), .O(n23827) );
  INV1S U14006 ( .I(n14056), .O(n14057) );
  INV2 U14007 ( .I(i_row[3]), .O(n23823) );
  INV2 U14008 ( .I(i_row[2]), .O(n14037) );
  NR2 U14009 ( .I1(n20892), .I2(n29455), .O(n20895) );
  AN4S U14010 ( .I1(n17542), .I2(n17541), .I3(n17540), .I4(n17539), .O(n17543)
         );
  AN4S U14011 ( .I1(n17705), .I2(n17704), .I3(n17703), .I4(n17702), .O(n17706)
         );
  MOAI1S U14012 ( .A1(n14914), .A2(n31371), .B1(n13837), .B2(img[763]), .O(
        n14872) );
  AN4S U14013 ( .I1(n17507), .I2(n17506), .I3(n17505), .I4(n17504), .O(n17508)
         );
  AN4S U14014 ( .I1(n17565), .I2(n17564), .I3(n17563), .I4(n17562), .O(n17566)
         );
  AN4S U14015 ( .I1(n19028), .I2(n19027), .I3(n19026), .I4(n19025), .O(n19029)
         );
  AN4S U14016 ( .I1(n18967), .I2(n18966), .I3(n18965), .I4(n18964), .O(n18968)
         );
  AN4S U14017 ( .I1(n18901), .I2(n18900), .I3(n18899), .I4(n18898), .O(n18902)
         );
  ND2 U14018 ( .I1(n16586), .I2(n16585), .O(n20559) );
  ND2 U14019 ( .I1(n16556), .I2(n16555), .O(n20557) );
  MOAI1S U14020 ( .A1(n15631), .A2(n31822), .B1(n13879), .B2(img[444]), .O(
        n15303) );
  MOAI1S U14021 ( .A1(n15631), .A2(n31906), .B1(n13879), .B2(img[428]), .O(
        n15181) );
  AN4S U14022 ( .I1(n18823), .I2(n18822), .I3(n18821), .I4(n18820), .O(n18830)
         );
  AN4S U14023 ( .I1(n18685), .I2(n18684), .I3(n18683), .I4(n18682), .O(n18691)
         );
  ND2 U14024 ( .I1(n17342), .I2(n17341), .O(n20481) );
  AN4S U14025 ( .I1(n16792), .I2(n16791), .I3(n16790), .I4(n16789), .O(n16793)
         );
  BUF2 U14026 ( .I(n19200), .O(n13855) );
  ND2 U14027 ( .I1(n16546), .I2(n16545), .O(n20542) );
  AN4S U14028 ( .I1(n18215), .I2(n18214), .I3(n18213), .I4(n18212), .O(n18216)
         );
  AOI22S U14029 ( .A1(n19342), .A2(img[811]), .B1(n17862), .B2(img[1451]), .O(
        n14779) );
  ND2 U14030 ( .I1(n18981), .I2(n18980), .O(n20085) );
  AN4S U14031 ( .I1(n18633), .I2(n18632), .I3(n18631), .I4(n18630), .O(n18639)
         );
  AN4S U14032 ( .I1(n18596), .I2(n18595), .I3(n18594), .I4(n18593), .O(n18597)
         );
  ND2 U14033 ( .I1(n17248), .I2(n17247), .O(n20477) );
  ND2 U14034 ( .I1(n19251), .I2(n19250), .O(n20244) );
  MOAI1S U14035 ( .A1(n16725), .A2(n17656), .B1(n16721), .B2(n20439), .O(
        n15153) );
  MOAI1S U14036 ( .A1(n16708), .A2(n13927), .B1(n16711), .B2(n14174), .O(
        n15147) );
  INV1S U14037 ( .I(n15652), .O(n15806) );
  MOAI1S U14038 ( .A1(n15780), .A2(n30214), .B1(n13885), .B2(img[815]), .O(
        n15650) );
  INV3 U14039 ( .I(n13856), .O(n13787) );
  INV3 U14040 ( .I(n13873), .O(n13874) );
  ND2 U14041 ( .I1(n17389), .I2(n17388), .O(n20484) );
  ND2 U14042 ( .I1(n16899), .I2(n16898), .O(n20442) );
  ND2 U14043 ( .I1(n16889), .I2(n16888), .O(n20454) );
  ND3S U14044 ( .I1(n14876), .I2(n14875), .I3(n14874), .O(n14883) );
  ND2 U14045 ( .I1(n19072), .I2(n19071), .O(n19987) );
  ND3S U14046 ( .I1(n15485), .I2(n15484), .I3(n15483), .O(n15486) );
  ND3S U14047 ( .I1(n15094), .I2(n15093), .I3(n15092), .O(n15101) );
  ND2 U14048 ( .I1(n18649), .I2(n18648), .O(n19745) );
  ND2 U14049 ( .I1(n18564), .I2(n18563), .O(n19747) );
  AN4S U14050 ( .I1(n15319), .I2(n15318), .I3(n15317), .I4(n15316), .O(n15326)
         );
  INV2 U14051 ( .I(n13849), .O(n14189) );
  ND3S U14052 ( .I1(n20337), .I2(n20336), .I3(n20335), .O(n20338) );
  AN4S U14053 ( .I1(n15683), .I2(n15682), .I3(n15681), .I4(n15680), .O(n15690)
         );
  ND3S U14054 ( .I1(n14124), .I2(n14123), .I3(n14122), .O(n14131) );
  BUF2 U14055 ( .I(n14909), .O(n18819) );
  MOAI1S U14056 ( .A1(n15780), .A2(n31688), .B1(n13884), .B2(img[864]), .O(
        n14583) );
  ND2 U14057 ( .I1(n16915), .I2(n16914), .O(n20441) );
  AN4S U14058 ( .I1(n17112), .I2(n17111), .I3(n17110), .I4(n17109), .O(n17113)
         );
  ND3S U14059 ( .I1(n14921), .I2(n14920), .I3(n14919), .O(n17671) );
  NR2 U14060 ( .I1(n14783), .I2(n14782), .O(n17655) );
  ND3S U14061 ( .I1(n15136), .I2(n15135), .I3(n15134), .O(n16729) );
  ND3S U14062 ( .I1(n14966), .I2(n14965), .I3(n14964), .O(n16705) );
  ND3 U14063 ( .I1(n15326), .I2(n15325), .I3(n15324), .O(n17936) );
  ND2 U14064 ( .I1(n18817), .I2(n18816), .O(n20365) );
  AN4S U14065 ( .I1(n19739), .I2(n19738), .I3(n19737), .I4(n19736), .O(n19740)
         );
  ND3 U14066 ( .I1(n20096), .I2(n20095), .I3(n20094), .O(n23180) );
  AN4S U14067 ( .I1(n18327), .I2(n18326), .I3(n18325), .I4(n18324), .O(n18328)
         );
  MOAI1S U14068 ( .A1(n17672), .A2(n15142), .B1(n17680), .B2(n13839), .O(
        n14936) );
  ND3S U14069 ( .I1(n15713), .I2(n15712), .I3(n15711), .O(n15720) );
  ND3S U14070 ( .I1(n14442), .I2(n14441), .I3(n14440), .O(n14449) );
  MOAI1S U14071 ( .A1(n17678), .A2(n13946), .B1(n17680), .B2(n13846), .O(
        n14871) );
  OAI12H U14072 ( .B1(n21422), .B2(n21421), .A1(n21420), .O(n21470) );
  ND3S U14073 ( .I1(n15785), .I2(n15784), .I3(n15783), .O(n16245) );
  INV1S U14074 ( .I(n20587), .O(n17418) );
  ND3S U14075 ( .I1(n14558), .I2(n14557), .I3(n14556), .O(n14565) );
  ND3S U14076 ( .I1(n16480), .I2(n16479), .I3(n16478), .O(n16498) );
  INV2 U14077 ( .I(n13766), .O(n13804) );
  ND2 U14078 ( .I1(n17104), .I2(n17103), .O(n21053) );
  INV1S U14079 ( .I(n21071), .O(n27891) );
  NR3 U14080 ( .I1(n15475), .I2(n15474), .I3(n15473), .O(n15578) );
  NR2T U14081 ( .I1(n13822), .I2(n19473), .O(n19603) );
  ND3S U14082 ( .I1(n14700), .I2(n14699), .I3(n14698), .O(n14706) );
  NR2 U14083 ( .I1(n15759), .I2(n15758), .O(n15818) );
  NR2 U14084 ( .I1(n14485), .I2(n14484), .O(n14486) );
  INV1S U14085 ( .I(n22058), .O(n22118) );
  ND3S U14086 ( .I1(n29971), .I2(n14006), .I3(n14005), .O(n14007) );
  INV1S U14087 ( .I(img_size[3]), .O(n23932) );
  MOAI1S U14088 ( .A1(n28573), .A2(n26037), .B1(n28571), .B2(n26036), .O(
        n26038) );
  OAI12HS U14089 ( .B1(n13995), .B2(n13994), .A1(n13993), .O(n23851) );
  OA112 U14090 ( .C1(n20855), .C2(n22918), .A1(n22917), .B1(n22916), .O(n13914) );
  INV1S U14091 ( .I(n22668), .O(n22730) );
  FA1S U14092 ( .A(n15900), .B(n15899), .CI(n15898), .CO(n15908), .S(n21772)
         );
  NR2 U14093 ( .I1(n14702), .I2(n14701), .O(n14703) );
  FA1S U14094 ( .A(n22341), .B(n22340), .CI(n22339), .CO(n22370), .S(n22367)
         );
  INV1S U14095 ( .I(n22417), .O(n22479) );
  INV1S U14096 ( .I(n21810), .O(n21871) );
  INV2 U14097 ( .I(n22061), .O(n22121) );
  INV1S U14098 ( .I(gray_avg[2]), .O(n23456) );
  NR2 U14099 ( .I1(n23932), .I2(n24034), .O(n24240) );
  NR2 U14100 ( .I1(n24515), .I2(n24692), .O(n24520) );
  BUF3 U14101 ( .I(n28415), .O(n13808) );
  NR2 U14102 ( .I1(n24708), .I2(n24692), .O(n24229) );
  BUF2 U14103 ( .I(n28415), .O(n28292) );
  ND2P U14104 ( .I1(n24240), .I2(img_size[1]), .O(n24495) );
  NR2P U14105 ( .I1(n23983), .I2(n24098), .O(n24515) );
  OAI112HS U14106 ( .C1(n13818), .C2(n19438), .A1(n18143), .B1(n22934), .O(
        n21398) );
  FA1S U14107 ( .A(n15597), .B(n15596), .CI(n15595), .CO(n15904), .S(n15841)
         );
  FA1S U14108 ( .A(n15953), .B(n15952), .CI(n15951), .CO(n15955), .S(n15995)
         );
  FA1S U14109 ( .A(n22357), .B(n22356), .CI(n22355), .CO(n22400), .S(n22393)
         );
  INV1S U14110 ( .I(c_s[1]), .O(n23565) );
  MOAI1S U14111 ( .A1(n23455), .A2(n23456), .B1(n23456), .B2(n23455), .O(
        n23463) );
  INV1S U14112 ( .I(c_s[2]), .O(n14029) );
  OAI12HS U14113 ( .B1(n24105), .B2(n24466), .A1(n24748), .O(n28598) );
  NR2 U14114 ( .I1(n24229), .I2(n24520), .O(n28864) );
  OAI12HS U14115 ( .B1(n24563), .B2(n24466), .A1(n24758), .O(n29033) );
  ND3S U14116 ( .I1(n25903), .I2(n25552), .I3(n25551), .O(n25553) );
  INV1S U14117 ( .I(n23122), .O(n23129) );
  INV1S U14118 ( .I(n22860), .O(n22867) );
  INV1S U14119 ( .I(n22670), .O(n22909) );
  OAI12HS U14120 ( .B1(n23380), .B2(n23330), .A1(n23329), .O(n23375) );
  FA1S U14121 ( .A(n15858), .B(n15857), .CI(n15856), .CO(n15918), .S(n21783)
         );
  INV1S U14122 ( .I(n22419), .O(n22651) );
  INV1S U14123 ( .I(n21994), .O(n22001) );
  INV1S U14124 ( .I(n22246), .O(n22253) );
  ND3S U14125 ( .I1(temp_cnt[2]), .I2(n29547), .I3(n29545), .O(n29544) );
  INV2 U14126 ( .I(in_valid2), .O(n29962) );
  ND2 U14127 ( .I1(n23587), .I2(n23561), .O(n30028) );
  ND3S U14128 ( .I1(n14032), .I2(n14011), .I3(n23694), .O(n30029) );
  INV2 U14129 ( .I(n13790), .O(n13854) );
  INV2 U14130 ( .I(n16799), .O(n13790) );
  INV3 U14131 ( .I(n14299), .O(n15315) );
  INV3 U14132 ( .I(n16468), .O(n17875) );
  BUF3 U14133 ( .I(n28318), .O(n28347) );
  INV1CK U14134 ( .I(n24700), .O(n28318) );
  OR2 U14135 ( .I1(n14146), .I2(n14213), .O(n13929) );
  MXL2HS U14136 ( .A(n21656), .B(n21655), .S(n21654), .OB(n13765) );
  MXL2HS U14137 ( .A(n29513), .B(n20385), .S(n21654), .OB(n21653) );
  INV1S U14138 ( .I(n23956), .O(n28043) );
  BUF1CK U14139 ( .I(n28043), .O(n28254) );
  BUF1CK U14140 ( .I(n28254), .O(n25444) );
  OR2 U14141 ( .I1(n14251), .I2(n14250), .O(n13766) );
  INV1S U14142 ( .I(n16186), .O(n23601) );
  BUF2 U14143 ( .I(n15652), .O(n13794) );
  BUF1S U14144 ( .I(n19245), .O(n16289) );
  BUF2 U14145 ( .I(n19245), .O(n13823) );
  BUF2 U14146 ( .I(n13842), .O(n19245) );
  BUF2 U14147 ( .I(n13842), .O(n15630) );
  BUF2 U14148 ( .I(n17885), .O(n20039) );
  INV6 U14149 ( .I(n13838), .O(n15800) );
  INV2 U14150 ( .I(n13872), .O(n13825) );
  INV1S U14151 ( .I(n13795), .O(n13831) );
  INV3 U14152 ( .I(n13840), .O(n15506) );
  NR2P U14153 ( .I1(n23623), .I2(n14047), .O(n16274) );
  INV1S U14154 ( .I(n13840), .O(n13795) );
  BUF1CK U14155 ( .I(n23918), .O(n24374) );
  BUF2 U14156 ( .I(n24193), .O(n25062) );
  BUF1CK U14157 ( .I(n24374), .O(n13779) );
  BUF1CK U14158 ( .I(n24193), .O(n13775) );
  BUF1CK U14159 ( .I(n23918), .O(n24193) );
  INV1S U14160 ( .I(n24699), .O(n23918) );
  BUF1CK U14161 ( .I(n23918), .O(n23941) );
  BUF1S U14162 ( .I(n29124), .O(n13899) );
  BUF1CK U14163 ( .I(n29258), .O(n13904) );
  BUF1S U14164 ( .I(n29124), .O(n29258) );
  BUF1CK U14165 ( .I(n29124), .O(n13819) );
  NR2T U14166 ( .I1(n23919), .I2(n24700), .O(n29124) );
  BUF1S U14167 ( .I(n29124), .O(n13902) );
  BUF1CK U14168 ( .I(n29124), .O(n13770) );
  BUF1S U14169 ( .I(n29124), .O(n13900) );
  BUF1S U14170 ( .I(n29124), .O(n13901) );
  BUF1CK U14171 ( .I(n29258), .O(n13905) );
  BUF1CK U14172 ( .I(n29258), .O(n13820) );
  MUX2S U14173 ( .A(n25640), .B(img[722]), .S(n29176), .O(n12810) );
  MUX2S U14174 ( .A(n25652), .B(img[746]), .S(n29112), .O(n12782) );
  MUX2S U14175 ( .A(n28243), .B(img[1064]), .S(n29115), .O(n12468) );
  MUX2S U14176 ( .A(n28202), .B(img[1712]), .S(n28722), .O(n11820) );
  MUX2S U14177 ( .A(n28233), .B(img[1576]), .S(n28729), .O(n11956) );
  MUX2S U14178 ( .A(n28238), .B(img[1552]), .S(n28736), .O(n11980) );
  MUX2S U14179 ( .A(n27545), .B(img[707]), .S(n28886), .O(n12825) );
  MUX2S U14180 ( .A(img[915]), .B(n27321), .S(n29061), .O(n12617) );
  MUX2S U14181 ( .A(n26927), .B(img[737]), .S(n29204), .O(n12795) );
  MUX2S U14182 ( .A(n28223), .B(img[1584]), .S(n28750), .O(n11948) );
  MUX2S U14183 ( .A(n27813), .B(img[731]), .S(n29377), .O(n12799) );
  MUX2S U14184 ( .A(n25759), .B(img[762]), .S(n29433), .O(n12766) );
  MUX2S U14185 ( .A(n25928), .B(img[730]), .S(n29377), .O(n12798) );
  MUX2S U14186 ( .A(img[1477]), .B(n26407), .S(n28872), .O(n12055) );
  MUX2S U14187 ( .A(img[1789]), .B(n26137), .S(n28941), .O(n11745) );
  ND3S U14188 ( .I1(n27769), .I2(n27393), .I3(n27392), .O(n27394) );
  ND3S U14189 ( .I1(n27769), .I2(n27410), .I3(n27409), .O(n27411) );
  BUF4 U14190 ( .I(n26583), .O(n13767) );
  BUF6 U14191 ( .I(n27769), .O(n13768) );
  BUF6CK U14192 ( .I(n25903), .O(n13769) );
  AOI12HP U14193 ( .B1(n28576), .B2(n28575), .A1(n28574), .O(n29278) );
  ND2 U14194 ( .I1(n21379), .I2(n21378), .O(n21381) );
  XNR2HS U14195 ( .I1(n21215), .I2(n21214), .O(n21207) );
  ND2S U14196 ( .I1(n23094), .I2(n23093), .O(n23120) );
  ND2S U14197 ( .I1(n22578), .I2(n22577), .O(n22597) );
  ND2 U14198 ( .I1(n24597), .I2(n24633), .O(n29481) );
  ND2 U14199 ( .I1(n24760), .I2(n24003), .O(n28666) );
  ND2 U14200 ( .I1(n24633), .I2(n24632), .O(n29380) );
  ND2S U14201 ( .I1(n22766), .I2(n22765), .O(n22870) );
  ND2 U14202 ( .I1(n24590), .I2(n24589), .O(n29142) );
  ND2 U14203 ( .I1(n24760), .I2(n24426), .O(n28889) );
  ND2 U14204 ( .I1(n24633), .I2(n24625), .O(n29374) );
  ND2 U14205 ( .I1(n24750), .I2(n24524), .O(n29106) );
  ND2 U14206 ( .I1(n24750), .I2(n24207), .O(n29230) );
  ND2 U14207 ( .I1(n24750), .I2(n24417), .O(n28883) );
  ND2 U14208 ( .I1(n24129), .I2(n23951), .O(n28620) );
  ND2 U14209 ( .I1(n24590), .I2(n24760), .O(n29173) );
  ND2 U14210 ( .I1(n24750), .I2(n24572), .O(n29170) );
  ND2 U14211 ( .I1(n24750), .I2(n24629), .O(n29371) );
  ND2 U14212 ( .I1(n24129), .I2(n24750), .O(n28659) );
  ND2 U14213 ( .I1(n24750), .I2(n24749), .O(n29427) );
  AO12 U14214 ( .B1(n24203), .B2(n24509), .A1(n24319), .O(n29255) );
  ND2 U14215 ( .I1(n24750), .I2(n24678), .O(n29328) );
  ND2 U14216 ( .I1(n24590), .I2(n24575), .O(n29166) );
  ND2 U14217 ( .I1(n24633), .I2(n24606), .O(n29348) );
  ND2 U14218 ( .I1(n24052), .I2(n24590), .O(n28701) );
  ND2 U14219 ( .I1(n24130), .I2(n24129), .O(n28792) );
  ND2 U14220 ( .I1(n24294), .I2(n24633), .O(n28951) );
  ND2 U14221 ( .I1(n24267), .I2(n24633), .O(n28922) );
  ND2 U14222 ( .I1(n24336), .I2(n24633), .O(n28993) );
  ND2 U14223 ( .I1(n24736), .I2(n24735), .O(n29416) );
  ND2 U14224 ( .I1(n24469), .I2(n24590), .O(n29047) );
  AO12 U14225 ( .B1(n24463), .B2(n24444), .A1(n24541), .O(n28818) );
  ND2 U14226 ( .I1(n24091), .I2(n24129), .O(n28750) );
  ND2 U14227 ( .I1(n24308), .I2(n24633), .O(n29185) );
  ND2 U14228 ( .I1(n24113), .I2(n24590), .O(n28771) );
  OR2S U14229 ( .I1(n22735), .I2(n22736), .O(n22895) );
  AO12 U14230 ( .B1(n24476), .B2(n24134), .A1(n24462), .O(n28617) );
  AO12 U14231 ( .B1(n24277), .B2(n24727), .A1(n24263), .O(n28941) );
  AO12 U14232 ( .B1(n24351), .B2(n24134), .A1(n24462), .O(n28796) );
  AO12 U14233 ( .B1(n24476), .B2(n24350), .A1(n24669), .O(n29240) );
  AO12 U14234 ( .B1(n24304), .B2(n24134), .A1(n24462), .O(n28754) );
  AO12 U14235 ( .B1(n24250), .B2(n24542), .A1(n24263), .O(n28683) );
  AO12 U14236 ( .B1(n24351), .B2(n24346), .A1(n24345), .O(n29004) );
  AO12 U14237 ( .B1(n24304), .B2(n24346), .A1(n24345), .O(n28962) );
  AO12 U14238 ( .B1(n24351), .B2(n24670), .A1(n24235), .O(n28789) );
  AO12 U14239 ( .B1(n24250), .B2(n24134), .A1(n24462), .O(n28698) );
  AO12 U14240 ( .B1(n24277), .B2(n24346), .A1(n24345), .O(n28933) );
  AO12 U14241 ( .B1(n24351), .B2(n24766), .A1(n24726), .O(n28785) );
  AO12 U14242 ( .B1(n24277), .B2(n24670), .A1(n24263), .O(n28719) );
  AO12 U14243 ( .B1(n24277), .B2(n24350), .A1(n24669), .O(n28929) );
  AO12 U14244 ( .B1(n24351), .B2(n24350), .A1(n24669), .O(n29000) );
  AO12 U14245 ( .B1(n24351), .B2(n24398), .A1(n24716), .O(n29018) );
  AO12 U14246 ( .B1(n24250), .B2(n24670), .A1(n24235), .O(n28690) );
  AO12 U14247 ( .B1(n24250), .B2(n24398), .A1(n24716), .O(n28919) );
  AO12 U14248 ( .B1(n24277), .B2(n24766), .A1(n24726), .O(n28715) );
  AO12 U14249 ( .B1(n24250), .B2(n24727), .A1(n24235), .O(n28911) );
  AO12 U14250 ( .B1(n24250), .B2(n24346), .A1(n24345), .O(n28903) );
  AN2S U14251 ( .I1(n27893), .I2(n21638), .O(n21307) );
  ND2 U14252 ( .I1(row[3]), .I2(n24012), .O(n23902) );
  HA1S U14253 ( .A(n15852), .B(n15851), .C(n15854), .S(n21788) );
  HA1S U14254 ( .A(n15836), .B(n15835), .C(n15889), .S(n15595) );
  INV2 U14255 ( .I(n22669), .O(n22776) );
  MOAI1H U14256 ( .A1(n21590), .A2(n21591), .B1(n21591), .B2(n21590), .O(
        n23438) );
  INV2 U14257 ( .I(n21805), .O(n13814) );
  INV3 U14258 ( .I(n21803), .O(n13812) );
  MXL2H U14259 ( .A(n20435), .B(n21336), .S(n20809), .OB(n29445) );
  ND3P U14260 ( .I1(n20377), .I2(n20376), .I3(n20375), .O(n22669) );
  OAI112HS U14261 ( .C1(n18318), .C2(n19235), .A1(n18317), .B1(n18316), .O(
        n22931) );
  ND2 U14262 ( .I1(n22915), .I2(n20809), .O(n19437) );
  ND3S U14263 ( .I1(n20306), .I2(n20305), .I3(n20304), .O(n20307) );
  INV2 U14264 ( .I(n18492), .O(n18489) );
  INV2 U14265 ( .I(n24665), .O(n24726) );
  AOI22S U14266 ( .A1(n19500), .A2(n20364), .B1(n20314), .B2(n19500), .O(
        n19502) );
  AOI22S U14267 ( .A1(n17957), .A2(n20371), .B1(n19533), .B2(n17957), .O(
        n17960) );
  AOI13HS U14268 ( .B1(n14939), .B2(n14938), .B3(n14937), .A1(n20969), .O(
        n19514) );
  ND2 U14269 ( .I1(n18483), .I2(n18482), .O(n18492) );
  ND2 U14270 ( .I1(n19532), .I2(n19531), .O(n19539) );
  NR3 U14271 ( .I1(n14931), .I2(n14930), .I3(n14929), .O(n14939) );
  ND2S U14272 ( .I1(n16225), .I2(n16224), .O(n16260) );
  ND2 U14273 ( .I1(n14013), .I2(c_s[2]), .O(n14032) );
  ND2 U14274 ( .I1(n16036), .I2(n16035), .O(n20619) );
  NR2 U14275 ( .I1(n14908), .I2(n14907), .O(n17672) );
  ND2 U14276 ( .I1(n18425), .I2(n18424), .O(n19834) );
  INV4 U14277 ( .I(n24722), .O(n24692) );
  ND3S U14278 ( .I1(n15610), .I2(n15609), .I3(n15608), .O(n15611) );
  AN4S U14279 ( .I1(n15269), .I2(n15268), .I3(n15267), .I4(n15266), .O(n15276)
         );
  ND2 U14280 ( .I1(n18994), .I2(n18993), .O(n20070) );
  AN4S U14281 ( .I1(n18689), .I2(n18688), .I3(n18687), .I4(n18686), .O(n18690)
         );
  AN4S U14282 ( .I1(n18710), .I2(n18709), .I3(n18708), .I4(n18707), .O(n18711)
         );
  AN4S U14283 ( .I1(n15805), .I2(n15804), .I3(n15803), .I4(n15802), .O(n15814)
         );
  AN4S U14284 ( .I1(n18828), .I2(n18827), .I3(n18826), .I4(n18825), .O(n18829)
         );
  AN4S U14285 ( .I1(n15725), .I2(n15724), .I3(n15723), .I4(n15722), .O(n15732)
         );
  AN4S U14286 ( .I1(n18627), .I2(n18626), .I3(n18625), .I4(n18624), .O(n18628)
         );
  ND3S U14287 ( .I1(n15737), .I2(n15736), .I3(n15735), .O(n15744) );
  BUF1 U14288 ( .I(n27746), .O(n13771) );
  BUF1 U14289 ( .I(n28382), .O(n13772) );
  BUF1 U14290 ( .I(n28840), .O(n13773) );
  INV2 U14291 ( .I(n29526), .O(n13774) );
  ND3 U14292 ( .I1(n15690), .I2(n15689), .I3(n15688), .O(n16244) );
  ND2 U14293 ( .I1(n18391), .I2(n18390), .O(n19825) );
  BUF1 U14294 ( .I(n29414), .O(n13776) );
  BUF1 U14295 ( .I(n28083), .O(n13777) );
  BUF1 U14296 ( .I(n27990), .O(n13778) );
  AN4S U14297 ( .I1(n17475), .I2(n17474), .I3(n17473), .I4(n17472), .O(n17476)
         );
  AN4S U14298 ( .I1(n15491), .I2(n15490), .I3(n15489), .I4(n15488), .O(n15498)
         );
  AN4S U14299 ( .I1(n18062), .I2(n18061), .I3(n18060), .I4(n18059), .O(n18063)
         );
  BUF1 U14300 ( .I(n26822), .O(n13780) );
  AN4S U14301 ( .I1(n15777), .I2(n15776), .I3(n15775), .I4(n15774), .O(n15785)
         );
  ND3S U14302 ( .I1(n14634), .I2(n14633), .I3(n14632), .O(n14641) );
  AN4S U14303 ( .I1(n18678), .I2(n18677), .I3(n18676), .I4(n18675), .O(n18679)
         );
  BUF3 U14304 ( .I(n23918), .O(n13781) );
  AN4S U14305 ( .I1(n18793), .I2(n18792), .I3(n18791), .I4(n18790), .O(n18794)
         );
  AN4S U14306 ( .I1(n18805), .I2(n18804), .I3(n18803), .I4(n18802), .O(n18806)
         );
  BUF3 U14307 ( .I(n28908), .O(n13782) );
  AN4S U14308 ( .I1(n17554), .I2(n17553), .I3(n17552), .I4(n17551), .O(n17555)
         );
  BUF3 U14309 ( .I(n18946), .O(n18935) );
  BUF2 U14310 ( .I(n18148), .O(n18988) );
  INV2 U14311 ( .I(n17828), .O(n13851) );
  BUF3 U14312 ( .I(n18946), .O(n19956) );
  BUF2 U14313 ( .I(n18148), .O(n19649) );
  NR2 U14314 ( .I1(n23797), .I2(n16172), .O(n16178) );
  INV3 U14315 ( .I(n13881), .O(n13882) );
  ND2 U14316 ( .I1(n13956), .I2(n13955), .O(n13958) );
  INV6 U14317 ( .I(n15801), .O(n13876) );
  INV4 U14318 ( .I(n17679), .O(n13830) );
  BUF2 U14319 ( .I(n15568), .O(n13784) );
  BUF4 U14320 ( .I(n19851), .O(n13859) );
  INV4 U14321 ( .I(n13872), .O(n13785) );
  BUF6 U14322 ( .I(n13828), .O(n13786) );
  BUF3 U14323 ( .I(n14909), .O(n20104) );
  BUF3 U14324 ( .I(n14909), .O(n18797) );
  BUF6 U14325 ( .I(n14189), .O(n13788) );
  BUF1 U14326 ( .I(n13945), .O(n17679) );
  INV12 U14327 ( .I(n14392), .O(n13789) );
  INV6 U14328 ( .I(n14044), .O(n15765) );
  BUF1 U14329 ( .I(n14044), .O(n17550) );
  BUF6 U14330 ( .I(n20103), .O(n13836) );
  BUF8CK U14331 ( .I(n17880), .O(n19710) );
  BUF3 U14332 ( .I(n14909), .O(n19411) );
  INV4 U14333 ( .I(n13927), .O(n13791) );
  BUF3 U14334 ( .I(n14909), .O(n19290) );
  BUF1 U14335 ( .I(n15561), .O(n13792) );
  BUF2 U14336 ( .I(n17418), .O(n13793) );
  BUF1 U14337 ( .I(n14044), .O(n13796) );
  BUF12CK U14338 ( .I(n16189), .O(n13797) );
  BUF1 U14339 ( .I(n13845), .O(n13799) );
  BUF8CK U14340 ( .I(n17880), .O(n13800) );
  BUF6 U14341 ( .I(n14555), .O(n13838) );
  BUF6 U14342 ( .I(n14909), .O(n13801) );
  AN2 U14343 ( .I1(n16170), .I2(n16169), .O(n16171) );
  ND2 U14344 ( .I1(n29969), .I2(n14029), .O(n23682) );
  ND2 U14345 ( .I1(n13989), .I2(act[11]), .O(n13990) );
  ND2S U14346 ( .I1(n13986), .I2(act[2]), .O(n13982) );
  ND2P U14347 ( .I1(n14050), .I2(n14056), .O(n16008) );
  BUF1 U14348 ( .I(n20039), .O(n13802) );
  INV12 U14349 ( .I(n15674), .O(n13803) );
  ND2 U14350 ( .I1(n13989), .I2(act[10]), .O(n13963) );
  NR2P U14351 ( .I1(act_ptr[2]), .I2(n13959), .O(n13987) );
  INV3 U14352 ( .I(n23623), .O(n14050) );
  INV2 U14353 ( .I(img_size[0]), .O(n28540) );
  INV2 U14354 ( .I(act_ptr[1]), .O(n13959) );
  BUF2 U14355 ( .I(img_size[2]), .O(n23900) );
  ND3 U14356 ( .I1(c_s[0]), .I2(c_s[1]), .I3(c_s[2]), .O(n29910) );
  BUF3 U14357 ( .I(rst_n), .O(n13805) );
  MUX2S U14358 ( .A(n23995), .B(img[823]), .S(n28659), .O(n12715) );
  MUX2S U14359 ( .A(n25872), .B(img[714]), .S(n28669), .O(n12814) );
  MUX2S U14360 ( .A(n25861), .B(img[818]), .S(n28659), .O(n12710) );
  MUX2S U14361 ( .A(img[476]), .B(n29365), .S(n29364), .O(n13056) );
  MUX2S U14362 ( .A(n26637), .B(img[733]), .S(n29377), .O(n12801) );
  MUX2S U14363 ( .A(n24761), .B(img[767]), .S(n29433), .O(n12771) );
  MUX2S U14364 ( .A(n26481), .B(img[717]), .S(n28669), .O(n12817) );
  MUX2S U14365 ( .A(n26462), .B(img[725]), .S(n29176), .O(n12807) );
  MUX2S U14366 ( .A(n26430), .B(img[709]), .S(n28886), .O(n12823) );
  MUX2S U14367 ( .A(n29335), .B(img[756]), .S(n29334), .O(n12776) );
  MUX2S U14368 ( .A(n26011), .B(img[706]), .S(n28886), .O(n12826) );
  MUX2S U14369 ( .A(n25976), .B(img[738]), .S(n29204), .O(n12794) );
  MUX2S U14370 ( .A(n24008), .B(img[719]), .S(n28669), .O(n12819) );
  MUX2S U14371 ( .A(img[468]), .B(n29164), .S(n29163), .O(n13064) );
  MUX2S U14372 ( .A(n25212), .B(img[718]), .S(n28669), .O(n12818) );
  MUX2S U14373 ( .A(n25205), .B(img[822]), .S(n28659), .O(n12714) );
  MUX2S U14374 ( .A(img[484]), .B(n29274), .S(n29273), .O(n13048) );
  MUX2S U14375 ( .A(img[900]), .B(n29396), .S(n29395), .O(n12632) );
  MUX2S U14376 ( .A(n25014), .B(img[758]), .S(n29334), .O(n12774) );
  MUX2S U14377 ( .A(img[499]), .B(n27682), .S(n29321), .O(n13033) );
  MUX2S U14378 ( .A(n25483), .B(img[754]), .S(n29334), .O(n12778) );
  MUX2S U14379 ( .A(n25390), .B(img[750]), .S(n29112), .O(n12786) );
  MUX2S U14380 ( .A(n25354), .B(img[726]), .S(n29176), .O(n12806) );
  MUX2S U14381 ( .A(n24857), .B(img[710]), .S(n28886), .O(n12822) );
  MUX2S U14382 ( .A(n29434), .B(img[764]), .S(n29433), .O(n12768) );
  MUX2S U14383 ( .A(n29378), .B(img[732]), .S(n29377), .O(n12800) );
  MUX2S U14384 ( .A(img[496]), .B(n28315), .S(n29321), .O(n13036) );
  MUX2S U14385 ( .A(n28335), .B(img[752]), .S(n29334), .O(n12780) );
  MUX2S U14386 ( .A(n28112), .B(img[760]), .S(n29433), .O(n12772) );
  MUX2S U14387 ( .A(img[896]), .B(n28091), .S(n29395), .O(n12636) );
  MUX2S U14388 ( .A(n28004), .B(img[704]), .S(n28886), .O(n12828) );
  MUX2S U14389 ( .A(n27887), .B(img[739]), .S(n29204), .O(n12793) );
  MUX2S U14390 ( .A(n27854), .B(img[763]), .S(n29433), .O(n12767) );
  MUX2S U14391 ( .A(n29177), .B(img[724]), .S(n29176), .O(n12808) );
  MUX2S U14392 ( .A(n27741), .B(img[715]), .S(n28669), .O(n12815) );
  MUX2S U14393 ( .A(n27703), .B(img[755]), .S(n29334), .O(n12777) );
  MUX2S U14394 ( .A(n29107), .B(img[876]), .S(n29106), .O(n12656) );
  MUX2S U14395 ( .A(n29113), .B(img[748]), .S(n29112), .O(n12784) );
  MUX2S U14396 ( .A(n28890), .B(img[700]), .S(n28889), .O(n12832) );
  MUX2S U14397 ( .A(n28884), .B(img[828]), .S(n28883), .O(n12704) );
  MUX2S U14398 ( .A(n28670), .B(img[716]), .S(n28669), .O(n12816) );
  MUX2S U14399 ( .A(n29208), .B(img[1188]), .S(n29207), .O(n12344) );
  MUX2S U14400 ( .A(n28526), .B(img[736]), .S(n29204), .O(n12796) );
  MUX2S U14401 ( .A(n28493), .B(img[712]), .S(n28669), .O(n12820) );
  MUX2S U14402 ( .A(n28486), .B(img[816]), .S(n28659), .O(n12716) );
  MUX2S U14403 ( .A(n24431), .B(img[711]), .S(n28886), .O(n12821) );
  MUX2S U14404 ( .A(n24580), .B(img[727]), .S(n29176), .O(n12805) );
  MUX2S U14405 ( .A(n28414), .B(img[728]), .S(n29377), .O(n12804) );
  MUX2S U14406 ( .A(n28379), .B(img[928]), .S(n29348), .O(n12604) );
  MUX2S U14407 ( .A(n29171), .B(img[852]), .S(n29170), .O(n12680) );
  MUX2S U14408 ( .A(n26993), .B(img[721]), .S(n29176), .O(n12811) );
  MUX2S U14409 ( .A(n26884), .B(img[729]), .S(n29377), .O(n12797) );
  MUX2S U14410 ( .A(n26731), .B(img[761]), .S(n29433), .O(n12765) );
  MUX2S U14411 ( .A(n27478), .B(img[723]), .S(n29176), .O(n12809) );
  MUX2S U14412 ( .A(n29428), .B(img[892]), .S(n29427), .O(n12640) );
  MUX2S U14413 ( .A(n27460), .B(img[939]), .S(n29142), .O(n12593) );
  MUX2S U14414 ( .A(n27350), .B(img[747]), .S(n29112), .O(n12783) );
  MUX2S U14415 ( .A(n27259), .B(img[745]), .S(n29112), .O(n12781) );
  MUX2S U14416 ( .A(n24687), .B(img[759]), .S(n29334), .O(n12773) );
  MUX2S U14417 ( .A(n29372), .B(img[860]), .S(n29371), .O(n12672) );
  MUX2S U14418 ( .A(n27226), .B(img[705]), .S(n28886), .O(n12827) );
  MUX2S U14419 ( .A(n27194), .B(img[713]), .S(n28669), .O(n12813) );
  MUX2S U14420 ( .A(n27188), .B(img[817]), .S(n28659), .O(n12709) );
  MUX2S U14421 ( .A(img[448]), .B(n27994), .S(n28857), .O(n13084) );
  MUX2S U14422 ( .A(img[450]), .B(n26000), .S(n28857), .O(n13082) );
  MUX2S U14423 ( .A(n28248), .B(img[1040]), .S(n29122), .O(n12492) );
  MUX2S U14424 ( .A(n28217), .B(img[1680]), .S(n28708), .O(n11852) );
  MUX2S U14425 ( .A(n28269), .B(img[1936]), .S(n28778), .O(n11596) );
  MUX2S U14426 ( .A(n28293), .B(img[1328]), .S(n28612), .O(n12204) );
  MUX2S U14427 ( .A(n28328), .B(img[1416]), .S(n28645), .O(n12116) );
  MUX2S U14428 ( .A(img[472]), .B(n28394), .S(n29364), .O(n13060) );
  MUX2S U14429 ( .A(img[498]), .B(n25463), .S(n29321), .O(n13034) );
  MUX2S U14430 ( .A(img[480]), .B(n28517), .S(n29273), .O(n13052) );
  MUX2S U14431 ( .A(n28274), .B(img[624]), .S(n29292), .O(n12908) );
  MUX2S U14432 ( .A(img[491]), .B(n27331), .S(n29084), .O(n13039) );
  MUX2S U14433 ( .A(img[483]), .B(n27878), .S(n29273), .O(n13049) );
  MUX2S U14434 ( .A(img[467]), .B(n27470), .S(n29163), .O(n13065) );
  MUX2S U14435 ( .A(n28080), .B(img[632]), .S(n29386), .O(n12900) );
  MUX2S U14436 ( .A(n28497), .B(img[608]), .S(n29286), .O(n12924) );
  MUX2S U14437 ( .A(img[1619]), .B(n27411), .S(n28733), .O(n11911) );
  MUX2S U14438 ( .A(img[1771]), .B(n27394), .S(n28712), .O(n11759) );
  MUX2S U14439 ( .A(img[1736]), .B(n28205), .S(n28726), .O(n11796) );
  MUX2S U14440 ( .A(img[1988]), .B(n29016), .S(n29015), .O(n11544) );
  MUX2S U14441 ( .A(img[1484]), .B(n28657), .S(n28656), .O(n12048) );
  MUX2S U14442 ( .A(img[1769]), .B(n27028), .S(n28712), .O(n11757) );
  MUX2S U14443 ( .A(img[1614]), .B(n25070), .S(n28754), .O(n11918) );
  MUX2S U14444 ( .A(img[1991]), .B(n24325), .S(n29015), .O(n11541) );
  MUX2S U14445 ( .A(img[1472]), .B(n27962), .S(n28872), .O(n12060) );
  MUX2S U14446 ( .A(img[2026]), .B(n25565), .S(n28782), .O(n11502) );
  MUX2S U14447 ( .A(img[1138]), .B(n25553), .S(n28761), .O(n12390) );
  ND3S U14448 ( .I1(n29278), .I2(n28655), .I3(n28654), .O(n28657) );
  ND3S U14449 ( .I1(n28415), .I2(n28204), .I3(n28203), .O(n28205) );
  ND3S U14450 ( .I1(n28415), .I2(n27961), .I3(n27960), .O(n27962) );
  INV4CK U14451 ( .I(n21458), .O(n21450) );
  ND3S U14452 ( .I1(n29278), .I2(n29014), .I3(n29013), .O(n29016) );
  BUF4 U14453 ( .I(n29278), .O(n13806) );
  BUF4 U14454 ( .I(n26583), .O(n13807) );
  INV1 U14455 ( .I(n21451), .O(n21384) );
  MUXB2 U14456 ( .EB(n21303), .A(n21302), .B(n21301), .S(n21300), .O(n21451)
         );
  ND2S U14457 ( .I1(n23379), .I2(n23378), .O(n23384) );
  AOI12HS U14458 ( .B1(n21909), .B2(n22006), .A1(n21908), .O(n21994) );
  ND2S U14459 ( .I1(n22245), .I2(n22244), .O(n22250) );
  ND2S U14460 ( .I1(n22257), .I2(n22256), .O(n22260) );
  ND2S U14461 ( .I1(n23128), .I2(n23127), .O(n23130) );
  ND2S U14462 ( .I1(n23139), .I2(n23138), .O(n23140) );
  ND2S U14463 ( .I1(n22621), .I2(n22620), .O(n22622) );
  ND2S U14464 ( .I1(n22603), .I2(n22602), .O(n22608) );
  ND2S U14465 ( .I1(n23374), .I2(n23369), .O(n23358) );
  ND2 U14466 ( .I1(n13909), .I2(n21476), .O(n21481) );
  ND2S U14467 ( .I1(n22263), .I2(n22262), .O(n22264) );
  INV1S U14468 ( .I(mult_x_431_n8), .O(n15913) );
  ND2S U14469 ( .I1(n21993), .I2(n21992), .O(n21998) );
  ND2S U14470 ( .I1(n22005), .I2(n22004), .O(n22008) );
  ND2S U14471 ( .I1(n23350), .I2(n23349), .O(n23373) );
  ND2S U14472 ( .I1(n22220), .I2(n22219), .O(n22239) );
  ND2 U14473 ( .I1(n24750), .I2(n24421), .O(n28879) );
  ND2S U14474 ( .I1(n21907), .I2(n21906), .O(n22004) );
  ND2 U14475 ( .I1(n24760), .I2(n24214), .O(n29204) );
  ND2 U14476 ( .I1(n24750), .I2(n23998), .O(n28663) );
  ND2 U14477 ( .I1(n24760), .I2(n24530), .O(n29112) );
  ND2 U14478 ( .I1(n24760), .I2(n24579), .O(n29176) );
  ND2 U14479 ( .I1(n24760), .I2(n24759), .O(n29433) );
  ND2 U14480 ( .I1(n24760), .I2(n24007), .O(n28669) );
  ND2 U14481 ( .I1(n24760), .I2(n24637), .O(n29377) );
  ND2 U14482 ( .I1(n24760), .I2(n24686), .O(n29334) );
  ND2 U14483 ( .I1(n24760), .I2(n24430), .O(n28886) );
  ND2S U14484 ( .I1(n22808), .I2(n22807), .O(n22858) );
  OR2S U14485 ( .I1(n23351), .I2(n23352), .O(n23369) );
  ND2P U14486 ( .I1(n24748), .I2(n24744), .O(n24750) );
  AO12 U14487 ( .B1(n24463), .B2(n24346), .A1(n24462), .O(n29218) );
  AO12 U14488 ( .B1(n24463), .B2(n24542), .A1(n24462), .O(n29044) );
  AO12 U14489 ( .B1(n24463), .B2(n24727), .A1(n24462), .O(n28814) );
  MOAI1 U14490 ( .A1(n21003), .A2(n21002), .B1(n22055), .B2(n21001), .O(n21005) );
  AO12 U14491 ( .B1(n24463), .B2(n24622), .A1(n24462), .O(n29211) );
  AO12 U14492 ( .B1(n24463), .B2(n24670), .A1(n24462), .O(n28595) );
  HA1S U14493 ( .A(n23204), .B(n23203), .C(n23211), .S(n23200) );
  HA1S U14494 ( .A(n23215), .B(n23214), .C(n23301), .S(n23219) );
  HA1S U14495 ( .A(n22994), .B(n22993), .C(n22987), .S(n23005) );
  HA1S U14496 ( .A(n22457), .B(n22456), .C(n22458), .S(n22468) );
  ND2 U14497 ( .I1(n23974), .I2(n23982), .O(n24664) );
  HA1S U14498 ( .A(n22471), .B(n22470), .C(n22464), .S(n22483) );
  INV3 U14499 ( .I(n23178), .O(n23292) );
  FA1S U14500 ( .A(n15891), .B(n15890), .CI(n15889), .CO(n21765), .S(n21768)
         );
  HA1S U14501 ( .A(n23232), .B(n23231), .C(n23228), .S(n23233) );
  FA1S U14502 ( .A(n15839), .B(n15838), .CI(n15837), .CO(n21767), .S(n15845)
         );
  HA1S U14503 ( .A(n22446), .B(n22445), .C(n22442), .S(n22492) );
  HA1S U14504 ( .A(n23193), .B(n23192), .C(n23194), .S(n23189) );
  HA1S U14505 ( .A(n22089), .B(n22088), .C(n22173), .S(n22093) );
  HA1S U14506 ( .A(n22120), .B(n22119), .C(n22115), .S(n22124) );
  FA1S U14507 ( .A(n15377), .B(n15376), .CI(n15375), .CO(n15844), .S(n15859)
         );
  FA1S U14508 ( .A(n15903), .B(n15902), .CI(n15901), .CO(n21771), .S(n21769)
         );
  HA1S U14509 ( .A(n22435), .B(n22434), .C(n22531), .S(n22430) );
  OR2P U14510 ( .I1(n23902), .I2(row[2]), .O(n24002) );
  HA1S U14511 ( .A(n22463), .B(n22462), .C(n22493), .S(n22496) );
  AN2S U14512 ( .I1(n17965), .I2(n21416), .O(n21417) );
  MOAI1 U14513 ( .A1(n28573), .A2(n25418), .B1(n28571), .B2(n25417), .O(n25419) );
  MOAI1 U14514 ( .A1(n28573), .A2(n23890), .B1(n28571), .B2(n23889), .O(n23891) );
  MOAI1 U14515 ( .A1(n28573), .A2(n24792), .B1(n28571), .B2(n24791), .O(n24793) );
  HA1S U14516 ( .A(n21870), .B(n21869), .C(n21866), .S(n22037) );
  HA1S U14517 ( .A(n22716), .B(n22715), .C(n22710), .S(n22717) );
  MOAI1 U14518 ( .A1(n28573), .A2(n26668), .B1(n28571), .B2(n26667), .O(n26669) );
  INV4CK U14519 ( .I(n22053), .O(n13809) );
  ND2S U14520 ( .I1(n21416), .I2(n20784), .O(n20785) );
  MOAI1 U14521 ( .A1(n28573), .A2(n28572), .B1(n28571), .B2(n28570), .O(n28574) );
  MOAI1 U14522 ( .A1(n28573), .A2(n27287), .B1(n28571), .B2(n27286), .O(n27288) );
  HA1S U14523 ( .A(n15877), .B(n15876), .C(n15893), .S(n15901) );
  HA1S U14524 ( .A(n22673), .B(n22672), .C(n22677), .S(n22743) );
  HA1S U14525 ( .A(n22687), .B(n22686), .C(n22694), .S(n22680) );
  HA1S U14526 ( .A(n15847), .B(n15846), .C(n15858), .S(n15853) );
  HA1S U14527 ( .A(n22698), .B(n22697), .C(n22781), .S(n22702) );
  HA1S U14528 ( .A(n21825), .B(n21824), .C(n21835), .S(n21826) );
  HA1S U14529 ( .A(n22709), .B(n22708), .C(n22674), .S(n22746) );
  INV2 U14530 ( .I(n22055), .O(n22168) );
  INV2 U14531 ( .I(n23186), .O(n23244) );
  OR2S U14532 ( .I1(n20784), .I2(n22054), .O(n20760) );
  NR2T U14533 ( .I1(n21330), .I2(n20499), .O(n29486) );
  INV2 U14534 ( .I(n23184), .O(n23299) );
  INV2 U14535 ( .I(n22062), .O(n13810) );
  INV4CK U14536 ( .I(n22411), .O(n13811) );
  INV2 U14537 ( .I(n23180), .O(n23295) );
  HA1S U14538 ( .A(n21839), .B(n21838), .C(n21921), .S(n21843) );
  HA1S U14539 ( .A(n21792), .B(n21791), .C(n21789), .S(PE_N49) );
  ND2P U14540 ( .I1(n22410), .I2(n20809), .O(n19461) );
  INV2 U14541 ( .I(n22662), .O(n22773) );
  OR2S U14542 ( .I1(n20776), .I2(n22418), .O(n20743) );
  INV2 U14543 ( .I(n29445), .O(n27263) );
  OR2S U14544 ( .I1(n20784), .I2(n23179), .O(n20700) );
  ND3P U14545 ( .I1(n13933), .I2(n16504), .I3(n16503), .O(n22054) );
  FA1S U14546 ( .A(n15884), .B(n15883), .CI(n15882), .CO(n15880), .S(n15909)
         );
  HA1S U14547 ( .A(n21690), .B(n21689), .C(n21697), .S(n22387) );
  OR2P U14548 ( .I1(n20168), .I2(n20167), .O(n23184) );
  INV1 U14549 ( .I(n26012), .O(n21596) );
  OR2S U14550 ( .I1(n20855), .I2(n22661), .O(n21125) );
  INV2 U14551 ( .I(n22661), .O(n22778) );
  ND3P U14552 ( .I1(n20302), .I2(n20301), .I3(n20300), .O(n22662) );
  AOI12HS U14553 ( .B1(n20298), .B2(n20363), .A1(n20297), .O(n20301) );
  HA1S U14554 ( .A(n23469), .B(n23468), .C(n23554), .S(PE_N65) );
  ND3P U14555 ( .I1(n20312), .I2(n20311), .I3(n20310), .O(n22663) );
  HA1S U14556 ( .A(n15984), .B(n15983), .C(n15982), .S(n21725) );
  INV2 U14557 ( .I(n21659), .O(n13813) );
  INV2 U14558 ( .I(n21658), .O(n22331) );
  HA1S U14559 ( .A(n15961), .B(n15960), .C(n15965), .S(n15962) );
  NR2 U14560 ( .I1(n19982), .I2(n13924), .O(n20009) );
  AOI12HS U14561 ( .B1(n20286), .B2(n20314), .A1(n20285), .O(n20289) );
  MXL2H U14562 ( .A(n20465), .B(n21333), .S(n20809), .OB(n26639) );
  INV2 U14563 ( .I(n29441), .O(n13815) );
  OR2 U14564 ( .I1(n14028), .I2(n23586), .O(n30027) );
  AOI22S U14565 ( .A1(n20372), .A2(n20364), .B1(n20363), .B2(n20372), .O(
        n20377) );
  INV4 U14566 ( .I(n21225), .O(n13818) );
  AOI13HS U14567 ( .B1(n15593), .B2(n15592), .B3(n15591), .A1(n20969), .O(
        n19474) );
  ND2S U14568 ( .I1(n16740), .I2(n19608), .O(n16691) );
  ND3S U14569 ( .I1(n20584), .I2(n20583), .I3(n20582), .O(n20600) );
  NR3 U14570 ( .I1(n15147), .I2(n15146), .I3(n15145), .O(n15156) );
  ND2 U14571 ( .I1(n18310), .I2(n18309), .O(n18315) );
  ND2 U14572 ( .I1(n19451), .I2(n19450), .O(n19457) );
  ND2P U14573 ( .I1(n17131), .I2(n17130), .O(n17191) );
  ND2S U14574 ( .I1(n20222), .I2(n20221), .O(n20228) );
  ND2S U14575 ( .I1(n20632), .I2(n20631), .O(n20633) );
  AN4S U14576 ( .I1(n16590), .I2(n16589), .I3(n16588), .I4(n16587), .O(n16667)
         );
  ND2S U14577 ( .I1(n20244), .I2(n20366), .O(n20226) );
  ND2 U14578 ( .I1(c_s[0]), .I2(n14021), .O(n14013) );
  BUF1 U14579 ( .I(n23941), .O(n29530) );
  BUF1 U14580 ( .I(n24193), .O(n29407) );
  ND2S U14581 ( .I1(n20244), .I2(n19818), .O(n20224) );
  BUF1 U14582 ( .I(n23941), .O(n24755) );
  ND2S U14583 ( .I1(n20585), .I2(n20580), .O(n16424) );
  BUF1 U14584 ( .I(n25062), .O(n28592) );
  BUF1 U14585 ( .I(n24193), .O(n29397) );
  ND2 U14586 ( .I1(n24612), .I2(n24694), .O(n24633) );
  BUF1 U14587 ( .I(n23941), .O(n28695) );
  ND2 U14588 ( .I1(n24758), .I2(n24563), .O(n24590) );
  NR2 U14589 ( .I1(n15413), .I2(n15412), .O(n16491) );
  ND2 U14590 ( .I1(n18447), .I2(n18446), .O(n19824) );
  BUF2 U14591 ( .I(n23941), .O(n28862) );
  ND2 U14592 ( .I1(n19325), .I2(n19324), .O(n20235) );
  BUF1 U14593 ( .I(n13781), .O(n29457) );
  ND2 U14594 ( .I1(n16849), .I2(n16848), .O(n20453) );
  ND3 U14595 ( .I1(n15814), .I2(n15813), .I3(n15812), .O(n16234) );
  BUF2 U14596 ( .I(n28043), .O(n28069) );
  NR2 U14597 ( .I1(n15612), .I2(n15611), .O(n16230) );
  BUF1 U14598 ( .I(n13781), .O(n28913) );
  BUF1 U14599 ( .I(n24374), .O(n27049) );
  AN2 U14600 ( .I1(n24240), .I2(n23973), .O(n23975) );
  ND3 U14601 ( .I1(n15703), .I2(n15702), .I3(n15701), .O(n16246) );
  ND2 U14602 ( .I1(n19355), .I2(n19354), .O(n20232) );
  AO12 U14603 ( .B1(n13781), .B2(n24035), .A1(n24345), .O(n24263) );
  ND2 U14604 ( .I1(n18371), .I2(n18370), .O(n19833) );
  ND2 U14605 ( .I1(n18917), .I2(n18916), .O(n20081) );
  BUF1 U14606 ( .I(n23941), .O(n25377) );
  ND2 U14607 ( .I1(n18415), .I2(n18414), .O(n19838) );
  INV2 U14608 ( .I(n24240), .O(n24694) );
  ND2 U14609 ( .I1(n16391), .I2(n16390), .O(n20594) );
  BUF1 U14610 ( .I(n28695), .O(n27511) );
  ND2 U14611 ( .I1(n19082), .I2(n19081), .O(n19997) );
  NR2 U14612 ( .I1(n15744), .I2(n15743), .O(n16241) );
  ND3 U14613 ( .I1(n15649), .I2(n15648), .I3(n15647), .O(n16236) );
  ND2 U14614 ( .I1(n19112), .I2(n19111), .O(n19996) );
  ND2 U14615 ( .I1(n19102), .I2(n19101), .O(n19995) );
  ND2 U14616 ( .I1(n19210), .I2(n19209), .O(n19986) );
  ND2 U14617 ( .I1(n18029), .I2(n18028), .O(n19882) );
  BUF2 U14618 ( .I(n24193), .O(n25591) );
  ND2 U14619 ( .I1(n18724), .I2(n18723), .O(n20151) );
  ND2 U14620 ( .I1(n18618), .I2(n18617), .O(n19744) );
  BUF1 U14621 ( .I(n29258), .O(n13903) );
  NR2 U14622 ( .I1(n15720), .I2(n15719), .O(n16239) );
  ND2 U14623 ( .I1(n19177), .I2(n19176), .O(n19989) );
  BUF2 U14624 ( .I(n28043), .O(n24313) );
  AN4S U14625 ( .I1(n17464), .I2(n17463), .I3(n17462), .I4(n17461), .O(n17465)
         );
  AN4S U14626 ( .I1(n15515), .I2(n15514), .I3(n15513), .I4(n15512), .O(n15522)
         );
  AN4S U14627 ( .I1(n17797), .I2(n17796), .I3(n17795), .I4(n17794), .O(n17798)
         );
  AN4S U14628 ( .I1(n16867), .I2(n16866), .I3(n16865), .I4(n16864), .O(n16868)
         );
  AN4S U14629 ( .I1(n15417), .I2(n15416), .I3(n15415), .I4(n15414), .O(n15424)
         );
  AN4S U14630 ( .I1(n17092), .I2(n17091), .I3(n17090), .I4(n17089), .O(n17093)
         );
  AN4S U14631 ( .I1(n16757), .I2(n16756), .I3(n16755), .I4(n16754), .O(n16764)
         );
  AN4S U14632 ( .I1(n15027), .I2(n15026), .I3(n15025), .I4(n15024), .O(n15034)
         );
  AN4S U14633 ( .I1(n17538), .I2(n17537), .I3(n17536), .I4(n17535), .O(n17544)
         );
  AN4S U14634 ( .I1(n18699), .I2(n18698), .I3(n18697), .I4(n18696), .O(n18700)
         );
  AN4S U14635 ( .I1(n15440), .I2(n15439), .I3(n15438), .I4(n15437), .O(n15447)
         );
  AN4S U14636 ( .I1(n14809), .I2(n14808), .I3(n14807), .I4(n14806), .O(n14816)
         );
  AN4S U14637 ( .I1(n16847), .I2(n16846), .I3(n16845), .I4(n16844), .O(n16848)
         );
  ND2 U14638 ( .I1(n16047), .I2(n16046), .O(n20609) );
  AN4S U14639 ( .I1(n17037), .I2(n17036), .I3(n17035), .I4(n17034), .O(n17038)
         );
  AN4S U14640 ( .I1(n18413), .I2(n18412), .I3(n18411), .I4(n18410), .O(n18414)
         );
  AN4S U14641 ( .I1(n17081), .I2(n17080), .I3(n17079), .I4(n17078), .O(n17082)
         );
  AN4S U14642 ( .I1(n19175), .I2(n19174), .I3(n19173), .I4(n19172), .O(n19176)
         );
  ND3 U14643 ( .I1(n24034), .I2(n24033), .I3(n24042), .O(n24345) );
  AN4S U14644 ( .I1(n16540), .I2(n16539), .I3(n16538), .I4(n16537), .O(n16546)
         );
  AN4S U14645 ( .I1(n18842), .I2(n18841), .I3(n18840), .I4(n18839), .O(n18843)
         );
  AN4S U14646 ( .I1(n16778), .I2(n16777), .I3(n16776), .I4(n16775), .O(n16784)
         );
  AN4S U14647 ( .I1(n14374), .I2(n14373), .I3(n14372), .I4(n14371), .O(n14381)
         );
  AN4S U14648 ( .I1(n17832), .I2(n17831), .I3(n17830), .I4(n17829), .O(n17833)
         );
  AN4S U14649 ( .I1(n16747), .I2(n16746), .I3(n16745), .I4(n16744), .O(n16753)
         );
  AN4S U14650 ( .I1(n17492), .I2(n17491), .I3(n17490), .I4(n17489), .O(n17498)
         );
  AN4S U14651 ( .I1(n16893), .I2(n16892), .I3(n16891), .I4(n16890), .O(n16899)
         );
  ND2 U14652 ( .I1(n18064), .I2(n18063), .O(n19896) );
  AN4S U14653 ( .I1(n17749), .I2(n17748), .I3(n17747), .I4(n17746), .O(n17750)
         );
  AN4S U14654 ( .I1(n15342), .I2(n15341), .I3(n15340), .I4(n15339), .O(n15350)
         );
  AN4S U14655 ( .I1(n16645), .I2(n16644), .I3(n16643), .I4(n16642), .O(n16651)
         );
  AN4S U14656 ( .I1(n18369), .I2(n18368), .I3(n18367), .I4(n18366), .O(n18370)
         );
  AN4S U14657 ( .I1(n16873), .I2(n16872), .I3(n16871), .I4(n16870), .O(n16879)
         );
  AN4S U14658 ( .I1(n17722), .I2(n17721), .I3(n17720), .I4(n17719), .O(n17728)
         );
  AN4S U14659 ( .I1(n17527), .I2(n17526), .I3(n17525), .I4(n17524), .O(n17533)
         );
  AN4S U14660 ( .I1(n14428), .I2(n14427), .I3(n14426), .I4(n14425), .O(n14435)
         );
  AN4S U14661 ( .I1(n17738), .I2(n17737), .I3(n17736), .I4(n17735), .O(n17739)
         );
  ND2 U14662 ( .I1(n19133), .I2(n19132), .O(n19998) );
  AN4S U14663 ( .I1(n16768), .I2(n16767), .I3(n16766), .I4(n16765), .O(n16774)
         );
  AN4S U14664 ( .I1(n19110), .I2(n19109), .I3(n19108), .I4(n19107), .O(n19111)
         );
  AN4S U14665 ( .I1(n18163), .I2(n18162), .I3(n18161), .I4(n18160), .O(n18164)
         );
  AN4S U14666 ( .I1(n17575), .I2(n17574), .I3(n17573), .I4(n17572), .O(n17576)
         );
  BUF1 U14667 ( .I(n28318), .O(n28083) );
  BUF1 U14668 ( .I(n28318), .O(n27746) );
  AN4S U14669 ( .I1(n18733), .I2(n18732), .I3(n18731), .I4(n18730), .O(n18734)
         );
  ND2 U14670 ( .I1(n23918), .I2(n23900), .O(n24034) );
  BUF1 U14671 ( .I(n28318), .O(n26822) );
  AN4S U14672 ( .I1(n17616), .I2(n17615), .I3(n17614), .I4(n17613), .O(n17623)
         );
  AN4S U14673 ( .I1(n18769), .I2(n18768), .I3(n18767), .I4(n18766), .O(n18770)
         );
  NR2 U14674 ( .I1(n15798), .I2(n15797), .O(n15828) );
  BUF1 U14675 ( .I(n28318), .O(n29414) );
  AN4S U14676 ( .I1(n17485), .I2(n17484), .I3(n17483), .I4(n17482), .O(n17486)
         );
  BUF1 U14677 ( .I(n28318), .O(n27990) );
  AN4S U14678 ( .I1(n17549), .I2(n17548), .I3(n17547), .I4(n17546), .O(n17556)
         );
  AN4S U14679 ( .I1(n16762), .I2(n16761), .I3(n16760), .I4(n16759), .O(n16763)
         );
  AN4S U14680 ( .I1(n16772), .I2(n16771), .I3(n16770), .I4(n16769), .O(n16773)
         );
  INV2 U14681 ( .I(n29526), .O(n13821) );
  AN4S U14682 ( .I1(n16508), .I2(n16507), .I3(n16506), .I4(n16505), .O(n16514)
         );
  AN4S U14683 ( .I1(n16987), .I2(n16986), .I3(n16985), .I4(n16984), .O(n16988)
         );
  AN4S U14684 ( .I1(n16993), .I2(n16992), .I3(n16991), .I4(n16990), .O(n16999)
         );
  AN4S U14685 ( .I1(n16833), .I2(n16832), .I3(n16831), .I4(n16830), .O(n16839)
         );
  AN4S U14686 ( .I1(n16997), .I2(n16996), .I3(n16995), .I4(n16994), .O(n16998)
         );
  ND2 U14687 ( .I1(n16370), .I2(n16369), .O(n20578) );
  AN4S U14688 ( .I1(n17027), .I2(n17026), .I3(n17025), .I4(n17024), .O(n17028)
         );
  AN4S U14689 ( .I1(n16857), .I2(n16856), .I3(n16855), .I4(n16854), .O(n16858)
         );
  AN4S U14690 ( .I1(n17716), .I2(n17715), .I3(n17714), .I4(n17713), .O(n17717)
         );
  AN4S U14691 ( .I1(n16883), .I2(n16882), .I3(n16881), .I4(n16880), .O(n16889)
         );
  NR2 U14692 ( .I1(n14641), .I2(n14640), .O(n17165) );
  BUF1 U14693 ( .I(n28318), .O(n28840) );
  AN4S U14694 ( .I1(n16594), .I2(n16593), .I3(n16592), .I4(n16591), .O(n16600)
         );
  ND2 U14695 ( .I1(n19122), .I2(n19121), .O(n20000) );
  AN4S U14696 ( .I1(n16278), .I2(n16277), .I3(n16276), .I4(n16275), .O(n16284)
         );
  AN4S U14697 ( .I1(n16803), .I2(n16802), .I3(n16801), .I4(n16800), .O(n16804)
         );
  BUF1 U14698 ( .I(n28318), .O(n28382) );
  ND2 U14699 ( .I1(n17073), .I2(n17072), .O(n21059) );
  AN4S U14700 ( .I1(n16809), .I2(n16808), .I3(n16807), .I4(n16806), .O(n16815)
         );
  AN4S U14701 ( .I1(n17057), .I2(n17056), .I3(n17055), .I4(n17054), .O(n17063)
         );
  ND2 U14702 ( .I1(n19188), .I2(n19187), .O(n19999) );
  AN4S U14703 ( .I1(n16813), .I2(n16812), .I3(n16811), .I4(n16810), .O(n16814)
         );
  INV1S U14704 ( .I(n13851), .O(n13852) );
  AN4S U14705 ( .I1(n18788), .I2(n18787), .I3(n18786), .I4(n18785), .O(n18795)
         );
  OR2 U14706 ( .I1(n23924), .I2(n24699), .O(n24033) );
  AN4S U14707 ( .I1(n16751), .I2(n16750), .I3(n16749), .I4(n16748), .O(n16752)
         );
  OR2 U14708 ( .I1(n14014), .I2(n30026), .O(n23561) );
  AN4S U14709 ( .I1(n17451), .I2(n17450), .I3(n17449), .I4(n17448), .O(n17452)
         );
  AN4S U14710 ( .I1(n18365), .I2(n18364), .I3(n18363), .I4(n18362), .O(n18371)
         );
  AN4S U14711 ( .I1(n18873), .I2(n18872), .I3(n18871), .I4(n18870), .O(n18879)
         );
  AN4S U14712 ( .I1(n17071), .I2(n17070), .I3(n17069), .I4(n17068), .O(n17072)
         );
  INV6 U14713 ( .I(n13851), .O(n13853) );
  AN4S U14714 ( .I1(n17007), .I2(n17006), .I3(n17005), .I4(n17004), .O(n17008)
         );
  AN4S U14715 ( .I1(n17017), .I2(n17016), .I3(n17015), .I4(n17014), .O(n17018)
         );
  OR2 U14716 ( .I1(n23897), .I2(n24700), .O(n23956) );
  AN4S U14717 ( .I1(n17531), .I2(n17530), .I3(n17529), .I4(n17528), .O(n17532)
         );
  BUF3 U14718 ( .I(n18946), .O(n19037) );
  BUF2 U14719 ( .I(n18148), .O(n20110) );
  INV6 U14720 ( .I(n13878), .O(n13879) );
  INV12 U14721 ( .I(n13911), .O(n13822) );
  ND3 U14722 ( .I1(n13996), .I2(n23895), .I3(n23851), .O(n23607) );
  ND3 U14723 ( .I1(n23854), .I2(n23853), .I3(n23852), .O(n23894) );
  BUF2 U14724 ( .I(n13795), .O(n13883) );
  INV2 U14725 ( .I(n13789), .O(n13824) );
  AN2 U14726 ( .I1(n24705), .I2(n23883), .O(n28571) );
  BUF1 U14727 ( .I(n15568), .O(n13826) );
  INV3 U14728 ( .I(n13790), .O(n13827) );
  INV1S U14729 ( .I(n18934), .O(n13868) );
  AO22S U14730 ( .A1(n23867), .A2(row[3]), .B1(n23757), .B2(n23756), .O(n23758) );
  INV2 U14731 ( .I(n18109), .O(n13828) );
  BUF1 U14732 ( .I(n14044), .O(n17561) );
  BUF3 U14733 ( .I(n13803), .O(n18773) );
  BUF1 U14734 ( .I(n13800), .O(n13829) );
  INV1 U14735 ( .I(n15113), .O(n19851) );
  INV4 U14736 ( .I(n14896), .O(n15799) );
  AN2 U14737 ( .I1(n24031), .I2(n23900), .O(n24025) );
  BUF2 U14738 ( .I(n14739), .O(n16353) );
  BUF3 U14739 ( .I(n13803), .O(n17864) );
  BUF3 U14740 ( .I(n13803), .O(n17816) );
  BUF1 U14741 ( .I(n14259), .O(n15448) );
  INV4 U14742 ( .I(n14896), .O(n19709) );
  NR2 U14743 ( .I1(n16176), .I2(n16175), .O(n16177) );
  BUF2 U14744 ( .I(n13886), .O(n16348) );
  ND3 U14745 ( .I1(n13965), .I2(n13964), .I3(n13963), .O(n13966) );
  ND3 U14746 ( .I1(n13971), .I2(n13970), .I3(n30031), .O(n13972) );
  ND3 U14747 ( .I1(n13976), .I2(n13975), .I3(act_ptr[0]), .O(n13977) );
  ND3 U14748 ( .I1(n23870), .I2(n23869), .I3(n23932), .O(n28544) );
  BUF1 U14749 ( .I(n14044), .O(n13832) );
  ND3 U14750 ( .I1(temp_cnt[1]), .I2(temp_cnt[2]), .I3(n29549), .O(n29550) );
  ND3 U14751 ( .I1(n23870), .I2(n23869), .I3(img_size[3]), .O(n26653) );
  BUF4 U14752 ( .I(n13803), .O(n13833) );
  ND3 U14753 ( .I1(n13982), .I2(n13981), .I3(act_ptr[0]), .O(n13995) );
  ND3 U14754 ( .I1(n13992), .I2(n13991), .I3(n13990), .O(n13993) );
  XNR2HS U14755 ( .I1(n23828), .I2(n23867), .O(n16172) );
  ND2 U14756 ( .I1(n23692), .I2(n23691), .O(n23693) );
  ND3 U14757 ( .I1(temp_cnt[1]), .I2(temp_cnt[2]), .I3(n29547), .O(n29548) );
  INV2 U14758 ( .I(n14266), .O(n15113) );
  ND3 U14759 ( .I1(temp_cnt[2]), .I2(n29549), .I3(n29545), .O(n29546) );
  ND3 U14760 ( .I1(temp_cnt[1]), .I2(n29549), .I3(n29542), .O(n29543) );
  ND2 U14761 ( .I1(n23897), .I2(n23919), .O(n23923) );
  BUF2 U14762 ( .I(n17418), .O(n13835) );
  ND3 U14763 ( .I1(temp_cnt[1]), .I2(n29547), .I3(n29542), .O(n29541) );
  BUF12CK U14764 ( .I(n16189), .O(n13837) );
  OR2 U14765 ( .I1(n23682), .I2(in_valid2), .O(n23652) );
  AN2 U14766 ( .I1(n24015), .I2(n24152), .O(n24134) );
  INV4 U14767 ( .I(n19462), .O(n13839) );
  OR2 U14768 ( .I1(n14012), .I2(c_s[1]), .O(N25894) );
  AN2 U14769 ( .I1(n24226), .I2(n24228), .O(n24444) );
  ND3 U14770 ( .I1(n23954), .I2(n23898), .I3(img_size[3]), .O(n23919) );
  INV4 U14771 ( .I(n16274), .O(n13840) );
  ND3 U14772 ( .I1(n23954), .I2(n13948), .I3(n23665), .O(n23897) );
  ND3 U14773 ( .I1(in_valid), .I2(n29552), .I3(n29551), .O(n29553) );
  INV3 U14774 ( .I(n16008), .O(n13842) );
  INV2 U14775 ( .I(n18196), .O(n13843) );
  ND2 U14776 ( .I1(n23690), .I2(n30004), .O(n23692) );
  BUF3 U14777 ( .I(n14258), .O(n13844) );
  ND2 U14778 ( .I1(n21501), .I2(c_s[0]), .O(n29968) );
  INV4 U14779 ( .I(n13947), .O(n13846) );
  AN2 U14780 ( .I1(n24019), .I2(n24152), .O(n24585) );
  OR2 U14781 ( .I1(row[3]), .I2(n24010), .O(n24098) );
  ND2 U14782 ( .I1(in_valid), .I2(n30025), .O(n30023) );
  INV4 U14783 ( .I(n13946), .O(n13847) );
  OR2 U14784 ( .I1(col[3]), .I2(col[2]), .O(n24234) );
  OR2 U14785 ( .I1(col[1]), .I2(col[0]), .O(n24233) );
  OR2 U14786 ( .I1(img_size[4]), .I2(img_size[5]), .O(n24698) );
  ND2 U14787 ( .I1(row[0]), .I2(row[1]), .O(n24099) );
  XNR2H U14788 ( .I1(img_size[0]), .I2(img_size[1]), .O(n23870) );
  OR2 U14789 ( .I1(row[1]), .I2(row[0]), .O(n24112) );
  ND3 U14790 ( .I1(n20348), .I2(n20347), .I3(n20346), .O(n20349) );
  NR3H U14791 ( .I1(n14603), .I2(n14602), .I3(n14601), .O(n14705) );
  AOI12HS U14792 ( .B1(n22599), .B2(n22598), .A1(n22594), .O(n22595) );
  ND3 U14793 ( .I1(n15012), .I2(n15011), .I3(n15010), .O(n16712) );
  AOI12H U14794 ( .B1(n21402), .B2(n21401), .A1(n21400), .O(n21406) );
  XNR2H U14795 ( .I1(n21473), .I2(n21472), .O(n21492) );
  XOR2HS U14796 ( .I1(n21471), .I2(n21470), .O(n21473) );
  ND2P U14797 ( .I1(n21344), .I2(n21343), .O(n21348) );
  XNR2H U14798 ( .I1(n21351), .I2(n21352), .O(n21369) );
  AOI22H U14799 ( .A1(n20373), .A2(n21117), .B1(n19625), .B2(n19818), .O(
        n17688) );
  FA1S U14800 ( .A(n15600), .B(n15599), .CI(n15598), .CO(n15840), .S(n15861)
         );
  NR2P U14801 ( .I1(n22475), .I2(n22528), .O(n22420) );
  XNR2HS U14802 ( .I1(n21207), .I2(n21216), .O(n21208) );
  OAI12HS U14803 ( .B1(n20957), .B2(n21596), .A1(n21081), .O(n20958) );
  XNR2HP U14804 ( .I1(n21285), .I2(n20992), .O(n21091) );
  ND3 U14805 ( .I1(n20985), .I2(n20984), .I3(n20983), .O(n20986) );
  NR2P U14806 ( .I1(n16498), .I2(n16497), .O(n20385) );
  AOI13H U14807 ( .B1(n29518), .B2(n29491), .B3(n29516), .A1(n29490), .O(
        n29495) );
  OAI112HS U14808 ( .C1(n29514), .C2(n29489), .A1(n29488), .B1(n29487), .O(
        n29490) );
  ND2P U14809 ( .I1(n16905), .I2(n16904), .O(n16966) );
  OAI12HS U14810 ( .B1(n22053), .B2(n21467), .A1(n17968), .O(n17969) );
  MXL2HS U14811 ( .A(mult_x_433_n6), .B(mult_x_433_n5), .S(mult_x_433_n9), 
        .OB(n22315) );
  INV1S U14812 ( .I(n21722), .O(n21703) );
  INV1 U14813 ( .I(n15652), .O(n14914) );
  AOI12HS U14814 ( .B1(n21989), .B2(n21988), .A1(n21984), .O(n21985) );
  INV1CK U14815 ( .I(n21804), .O(n21918) );
  ND3P U14816 ( .I1(n16451), .I2(n16450), .I3(n16452), .O(n21804) );
  INV1S U14817 ( .I(n17174), .O(n14715) );
  AOI112HS U14818 ( .C1(n18492), .C2(n20371), .A1(n18491), .B1(n18490), .O(
        n22940) );
  AOI12HP U14819 ( .B1(n25420), .B2(n28575), .A1(n25419), .O(n25903) );
  XNR2HP U14820 ( .I1(n21353), .I2(n21349), .O(n21352) );
  OAI12HP U14821 ( .B1(n21236), .B2(n21467), .A1(n20640), .O(n21353) );
  INV2 U14822 ( .I(n20644), .O(n29483) );
  OAI112H U14823 ( .C1(n18665), .C2(n19661), .A1(n18664), .B1(n18663), .O(
        n22926) );
  INV1CK U14824 ( .I(n21236), .O(n21238) );
  MOAI1 U14825 ( .A1(n16948), .A2(n15142), .B1(n16947), .B2(n13847), .O(n16949) );
  AOI12H U14826 ( .B1(n16965), .B2(n19533), .A1(n16964), .O(n16968) );
  OAI12H U14827 ( .B1(n22053), .B2(n20855), .A1(n21257), .O(n21258) );
  INV1CK U14828 ( .I(n21200), .O(n21128) );
  ND2 U14829 ( .I1(n24466), .I2(n24694), .O(n24148) );
  OR2T U14830 ( .I1(n24705), .I2(n28575), .O(n13908) );
  INV1S U14831 ( .I(n21452), .O(n21455) );
  OAI12H U14832 ( .B1(n29443), .B2(n27263), .A1(n21077), .O(n21078) );
  NR2P U14833 ( .I1(n17685), .I2(n17684), .O(n20679) );
  NR2 U14834 ( .I1(n22293), .I2(n13809), .O(n22072) );
  ND3 U14835 ( .I1(n16258), .I2(n16257), .I3(n16256), .O(n16259) );
  ND3HT U14836 ( .I1(n15819), .I2(n15818), .I3(n15817), .O(n21259) );
  MXL2H U14837 ( .A(n23187), .B(n20976), .S(n13822), .OB(n21071) );
  MOAI1 U14838 ( .A1(n17161), .A2(n13947), .B1(n17160), .B2(n20263), .O(n17162) );
  INV3 U14839 ( .I(n14896), .O(n15691) );
  OAI12HS U14840 ( .B1(n21102), .B2(n21101), .A1(n21100), .O(n21453) );
  MAO222 U14841 ( .A1(n21099), .B1(n23841), .C1(n21106), .O(n21100) );
  OAI112HS U14842 ( .C1(n21072), .C2(n22417), .A1(n20842), .B1(n22419), .O(
        n20843) );
  OAI12H U14843 ( .B1(n21391), .B2(n21085), .A1(n20854), .O(n20991) );
  OAI22S U14844 ( .A1(n29441), .A2(n21079), .B1(n21076), .B2(n29493), .O(
        n20695) );
  ND3 U14845 ( .I1(n20702), .I2(n20701), .I3(n20700), .O(n20703) );
  NR2F U14846 ( .I1(n21219), .I2(n21218), .O(n21456) );
  ND2T U14847 ( .I1(n21209), .I2(n21208), .O(n21219) );
  ND2P U14848 ( .I1(n19572), .I2(n19571), .O(n19580) );
  AOI22H U14849 ( .A1(n13892), .A2(img[987]), .B1(n19642), .B2(img[219]), .O(
        n14761) );
  OAI12H U14850 ( .B1(n23122), .B2(n23110), .A1(n23109), .O(n23117) );
  AOI12H U14851 ( .B1(n22930), .B2(n22932), .A1(n22931), .O(n13912) );
  OR2 U14852 ( .I1(n21288), .I2(n21287), .O(n21298) );
  OAI112HS U14853 ( .C1(n21805), .C2(n19494), .A1(n20653), .B1(n20652), .O(
        n20655) );
  OAI12HS U14854 ( .B1(n21595), .B2(n21245), .A1(n20651), .O(n20653) );
  ND2 U14855 ( .I1(n17628), .I2(n17638), .O(n17653) );
  INV1 U14856 ( .I(n20872), .O(n20916) );
  AOI12HS U14857 ( .B1(n19539), .B2(n19608), .A1(n19538), .O(n19540) );
  NR2 U14858 ( .I1(n15913), .I2(mult_x_431_n11), .O(n15914) );
  NR2P U14859 ( .I1(n15868), .I2(n21726), .O(n15887) );
  INV1CK U14860 ( .I(n20537), .O(n21726) );
  OAI12H U14861 ( .B1(n23508), .B2(n18134), .A1(n15157), .O(n20537) );
  OAI12H U14862 ( .B1(n22604), .B2(n22592), .A1(n22591), .O(n22599) );
  INV4CK U14863 ( .I(n22412), .O(n22528) );
  AOI12H U14864 ( .B1(n19908), .B2(n20363), .A1(n19907), .O(n19909) );
  INV1S U14865 ( .I(n17405), .O(n17406) );
  AOI22H U14866 ( .A1(n20358), .A2(n20063), .B1(n19818), .B2(n19903), .O(
        n19904) );
  OAI12HP U14867 ( .B1(n23848), .B2(n23846), .A1(n21089), .O(n21357) );
  BUF2 U14868 ( .I(n15568), .O(n19376) );
  NR2T U14869 ( .I1(n20673), .I2(n20672), .O(n21446) );
  OAI12HP U14870 ( .B1(n13816), .B2(n19438), .A1(n18319), .O(n29455) );
  INV2 U14871 ( .I(n20503), .O(n29442) );
  AOI12H U14872 ( .B1(n28534), .B2(n23848), .A1(n23847), .O(n23849) );
  BUF6 U14873 ( .I(n15356), .O(n20863) );
  NR2F U14874 ( .I1(n21091), .I2(n21092), .O(n21104) );
  BUF8CK U14875 ( .I(n17454), .O(n22932) );
  AOI12H U14876 ( .B1(n18662), .B2(n20373), .A1(n18661), .O(n18663) );
  ND2S U14877 ( .I1(n18660), .I2(n18659), .O(n18661) );
  ND2P U14878 ( .I1(n18655), .I2(n18654), .O(n18662) );
  AOI12HP U14879 ( .B1(n27289), .B2(n28575), .A1(n27288), .O(n27769) );
  AOI12H U14880 ( .B1(n21419), .B2(n21418), .A1(n21417), .O(n21422) );
  INV3 U14881 ( .I(n18718), .O(n13888) );
  ND2 U14882 ( .I1(n21202), .I2(n21156), .O(n21212) );
  MOAI1H U14883 ( .A1(n20821), .A2(n20820), .B1(n21596), .B2(n20903), .O(
        n20823) );
  MOAI1 U14884 ( .A1(n15698), .A2(n31788), .B1(n20038), .B2(img[1900]), .O(
        n15323) );
  MOAI1 U14885 ( .A1(n17937), .A2(n20421), .B1(n17936), .B2(n13846), .O(n17942) );
  OAI12H U14886 ( .B1(n20383), .B2(n21449), .A1(n17969), .O(n21393) );
  NR3 U14887 ( .I1(n15056), .I2(n15055), .I3(n15054), .O(n15063) );
  INV2 U14888 ( .I(n21081), .O(n26015) );
  XNR2H U14889 ( .I1(n21201), .I2(n21200), .O(n21215) );
  ND3 U14890 ( .I1(n15558), .I2(n15557), .I3(n15556), .O(n15559) );
  MUXB2 U14891 ( .EB(n20935), .A(n20934), .B(n20933), .S(n20932), .O(n21388)
         );
  AOI22S U14892 ( .A1(n29492), .A2(n29483), .B1(n19587), .B2(n19586), .O(
        n19588) );
  AOI12H U14893 ( .B1(n20912), .B2(n20911), .A1(n20910), .O(n21479) );
  FA1 U14894 ( .A(n23324), .B(n23323), .CI(n23322), .CO(n23328), .S(n23326) );
  ND3 U14895 ( .I1(n20226), .I2(n20225), .I3(n20224), .O(n20227) );
  NR2T U14896 ( .I1(n16255), .I2(n20691), .O(n21669) );
  MOAI1S U14897 ( .A1(n15780), .A2(n30121), .B1(n13885), .B2(img[807]), .O(
        n15686) );
  ND2T U14898 ( .I1(n21259), .I2(n20809), .O(n20855) );
  MUX2 U14899 ( .A(img[1203]), .B(n27650), .S(n28598), .O(n12329) );
  ND2 U14900 ( .I1(n21213), .I2(n21212), .O(n21217) );
  INV2 U14901 ( .I(i_col[2]), .O(n23792) );
  INV3 U14902 ( .I(n23846), .O(n21460) );
  AO12 U14903 ( .B1(n20637), .B2(n20636), .A1(n21346), .O(n23846) );
  NR2 U14904 ( .I1(n15986), .I2(n23525), .O(n15928) );
  FA1 U14905 ( .A(n21941), .B(n21940), .CI(n21939), .CO(n21963), .S(n21907) );
  OAI22S U14906 ( .A1(n21088), .A2(n29508), .B1(n21079), .B2(n29444), .O(
        n20961) );
  INV3 U14907 ( .I(n21228), .O(n21336) );
  OAI12H U14908 ( .B1(n29448), .B2(n13844), .A1(n14940), .O(n21228) );
  INV4CK U14909 ( .I(n16009), .O(n15652) );
  ND2T U14910 ( .I1(n22932), .I2(n20809), .O(n29448) );
  OAI12HS U14911 ( .B1(n22628), .B2(n22624), .A1(n22625), .O(n22616) );
  INV2 U14912 ( .I(n18297), .O(n18885) );
  MUX2 U14913 ( .A(mult_x_433_n11), .B(mult_x_433_n10), .S(mult_x_433_n14), 
        .O(mult_x_433_n9) );
  FA1 U14914 ( .A(n22393), .B(n22392), .CI(n22391), .CO(n22401), .S(
        mult_x_433_n42) );
  FA1S U14915 ( .A(n22363), .B(n22362), .CI(n22361), .CO(n22398), .S(n22391)
         );
  OAI12H U14916 ( .B1(n21457), .B2(n21085), .A1(n20989), .O(n20990) );
  XNR2H U14917 ( .I1(n21199), .I2(n20991), .O(n20992) );
  ND2 U14918 ( .I1(n18217), .I2(n18216), .O(n19677) );
  OAI12HP U14919 ( .B1(n19708), .B2(n19707), .A1(n20942), .O(n21079) );
  OR2T U14920 ( .I1(n13822), .I2(n23185), .O(n20942) );
  INV3CK U14921 ( .I(n16009), .O(n14044) );
  XNR2HP U14922 ( .I1(n21476), .I2(n21436), .O(n21349) );
  OAI112HS U14923 ( .C1(n21613), .C2(n21407), .A1(n21342), .B1(n21341), .O(
        n21344) );
  OAI12HS U14924 ( .B1(n21618), .B2(n28531), .A1(n21339), .O(n21342) );
  ND3 U14925 ( .I1(n14794), .I2(n14793), .I3(n14792), .O(n17654) );
  OAI12H U14926 ( .B1(n28536), .B2(n27893), .A1(n27892), .O(n27916) );
  ND3HT U14927 ( .I1(n21498), .I2(n21497), .I3(n21496), .O(n28536) );
  AOI12H U14928 ( .B1(n28534), .B2(n27891), .A1(n27890), .O(n27892) );
  AOI12HP U14929 ( .B1(n27916), .B2(n28575), .A1(n27915), .O(n28415) );
  AOI22HP U14930 ( .A1(n23848), .A2(n21449), .B1(n21009), .B2(n21008), .O(
        n21425) );
  ND2P U14931 ( .I1(n19741), .I2(n19740), .O(n20329) );
  BUF3 U14932 ( .I(n15568), .O(n19288) );
  OAI12H U14933 ( .B1(n21754), .B2(n21753), .A1(n21752), .O(n21761) );
  OAI12H U14934 ( .B1(n21751), .B2(n21750), .A1(n21749), .O(n21752) );
  INV2 U14935 ( .I(n21221), .O(n21799) );
  OAI12H U14936 ( .B1(n22942), .B2(n18134), .A1(n18484), .O(n21221) );
  ND2P U14937 ( .I1(n17283), .I2(n17282), .O(n20480) );
  AOI22H U14938 ( .A1(n21237), .A2(n13812), .B1(n20655), .B2(n20654), .O(
        n21280) );
  NR2P U14939 ( .I1(n20808), .I2(n20807), .O(n21386) );
  MXL2H U14940 ( .A(n29467), .B(n20674), .S(n21654), .OB(n21658) );
  XNR2HS U14941 ( .I1(n21363), .I2(n21375), .O(n21364) );
  AOI22S U14942 ( .A1(n29502), .A2(n29493), .B1(n29521), .B2(n29492), .O(
        n29494) );
  ND3 U14943 ( .I1(n19906), .I2(n19905), .I3(n19904), .O(n19907) );
  MOAI1 U14944 ( .A1(n17414), .A2(n13927), .B1(n17413), .B2(n13846), .O(n17415) );
  ND3 U14945 ( .I1(n14435), .I2(n14434), .I3(n14433), .O(n17413) );
  INV2 U14946 ( .I(n15113), .O(n18262) );
  AOI22H U14947 ( .A1(n21612), .A2(n20899), .B1(n20819), .B2(n20818), .O(
        n20821) );
  OAI12HP U14948 ( .B1(n19461), .B2(n22661), .A1(n20826), .O(n21200) );
  XOR2H U14949 ( .I1(n21217), .I2(n23844), .O(n21218) );
  ND2S U14950 ( .I1(n29510), .I2(n29464), .O(n29465) );
  ND2P U14951 ( .I1(n20160), .I2(n20159), .O(n20372) );
  OAI12HP U14952 ( .B1(n23845), .B2(n23848), .A1(n20990), .O(n21199) );
  BUF1 U14953 ( .I(n16002), .O(n13849) );
  BUF6 U14954 ( .I(n16002), .O(n13850) );
  ND2P U14955 ( .I1(n14050), .I2(n14054), .O(n16002) );
  INV3 U14956 ( .I(n14174), .O(n15142) );
  INV1S U14957 ( .I(n14896), .O(n19200) );
  OR2P U14958 ( .I1(n14250), .I2(n14213), .O(n13945) );
  INV1 U14959 ( .I(n15561), .O(n13856) );
  INV8 U14960 ( .I(n13857), .O(n13858) );
  INV1S U14961 ( .I(n14896), .O(n20191) );
  BUF6 U14962 ( .I(n16289), .O(n19193) );
  BUF1 U14963 ( .I(n19127), .O(n13860) );
  BUF3 U14964 ( .I(n19127), .O(n13861) );
  ND2P U14965 ( .I1(n23834), .I2(n14145), .O(n16468) );
  INV8 U14966 ( .I(n13838), .O(n15561) );
  INV4 U14967 ( .I(n16431), .O(n18109) );
  INV1S U14968 ( .I(n16064), .O(n13862) );
  INV2 U14969 ( .I(n13862), .O(n13863) );
  INV12 U14970 ( .I(n13848), .O(n14505) );
  BUF12CK U14971 ( .I(n14505), .O(n14822) );
  BUF12CK U14972 ( .I(n14822), .O(n18148) );
  BUF6CK U14973 ( .I(n18148), .O(n17810) );
  BUF3 U14974 ( .I(n17810), .O(n16037) );
  INV1S U14975 ( .I(n19318), .O(n13864) );
  INV2 U14976 ( .I(n13864), .O(n13865) );
  INV1S U14977 ( .I(n17779), .O(n13866) );
  INV3 U14978 ( .I(n13866), .O(n13867) );
  INV3 U14979 ( .I(n20855), .O(n21237) );
  INV1S U14980 ( .I(n13868), .O(n13869) );
  INV2 U14981 ( .I(n13868), .O(n13870) );
  INV3 U14982 ( .I(n13840), .O(n13871) );
  INV6CK U14983 ( .I(n13871), .O(n13872) );
  BUF6 U14984 ( .I(n19245), .O(n17382) );
  MOAI1S U14985 ( .A1(n15780), .A2(n30123), .B1(n13885), .B2(img[871]), .O(
        n15728) );
  NR3H U14986 ( .I1(n15708), .I2(n15707), .I3(n15706), .O(n15819) );
  BUF6 U14987 ( .I(n16353), .O(n17862) );
  BUF3 U14988 ( .I(n17886), .O(n17515) );
  INV6 U14989 ( .I(n15674), .O(n14909) );
  BUF3 U14990 ( .I(n13803), .O(n17793) );
  BUF3 U14991 ( .I(n13803), .O(n18983) );
  BUF3 U14992 ( .I(n13803), .O(n18958) );
  BUF3 U14993 ( .I(n13803), .O(n17335) );
  BUF3 U14994 ( .I(n19403), .O(n13877) );
  INV2 U14995 ( .I(n13834), .O(n13878) );
  BUF4 U14996 ( .I(n19258), .O(n13880) );
  INV6 U14997 ( .I(n14266), .O(n14896) );
  MOAI1 U14998 ( .A1(n15113), .A2(n30213), .B1(n15786), .B2(img[279]), .O(
        n15710) );
  MOAI1 U14999 ( .A1(n15113), .A2(n30263), .B1(n15786), .B2(img[271]), .O(
        n15734) );
  INV2 U15000 ( .I(n15721), .O(n13881) );
  INV3CK U15001 ( .I(n15653), .O(n16516) );
  AN4 U15002 ( .I1(n17053), .I2(n17052), .I3(n17051), .I4(n17050), .O(n17131)
         );
  INV6 U15003 ( .I(n13888), .O(n13890) );
  AN2T U15004 ( .I1(n14055), .I2(n14054), .O(n13931) );
  INV12 U15005 ( .I(n13891), .O(n13893) );
  NR2P U15006 ( .I1(n14047), .I2(n14058), .O(n18155) );
  BUF6 U15007 ( .I(n14286), .O(n13887) );
  INV2 U15008 ( .I(n13888), .O(n13889) );
  INV6CK U15009 ( .I(n17115), .O(n13891) );
  INV6 U15010 ( .I(n13891), .O(n13892) );
  INV6CK U15011 ( .I(n13834), .O(n13894) );
  INV2 U15012 ( .I(n13894), .O(n13895) );
  INV6 U15013 ( .I(n13894), .O(n13896) );
  AN2T U15014 ( .I1(n19700), .I2(n18142), .O(n20063) );
  ND2S U15015 ( .I1(n20863), .I2(n18142), .O(n20367) );
  ND2 U15016 ( .I1(n19495), .I2(n18142), .O(n19050) );
  ND2 U15017 ( .I1(n20345), .I2(n18142), .O(n20346) );
  NR2P U15018 ( .I1(n18141), .I2(n13822), .O(n18142) );
  BUF3 U15019 ( .I(n28529), .O(n13897) );
  BUF6 U15020 ( .I(n16016), .O(n17522) );
  BUF6 U15021 ( .I(n16189), .O(n13898) );
  NR2P U15022 ( .I1(n14047), .I2(n14046), .O(n16189) );
  NR2P U15023 ( .I1(n24766), .I2(n24726), .O(n24682) );
  INV6CK U15024 ( .I(n18109), .O(n19215) );
  INV6CK U15025 ( .I(n18297), .O(n19036) );
  INV12 U15026 ( .I(n14034), .O(n15786) );
  OA12 U15027 ( .B1(n23929), .B2(n23928), .A1(n24510), .O(n24462) );
  FA1S U15028 ( .A(rgb_value[15]), .B(rgb_value[7]), .CI(rgb_value[23]), .CO(
        n21527), .S(n21522) );
  AN2S U15029 ( .I1(n21416), .I2(n24769), .O(n21321) );
  OR2S U15030 ( .I1(n22324), .I2(n20948), .O(n20701) );
  ND2S U15031 ( .I1(n14133), .I2(n14132), .O(n16059) );
  ND2S U15032 ( .I1(n17430), .I2(n17429), .O(n17431) );
  ND2S U15033 ( .I1(img_size[3]), .I2(n23900), .O(n23857) );
  ND2S U15034 ( .I1(n23855), .I2(img_size[3]), .O(n23856) );
  OR2S U15035 ( .I1(n23900), .I2(img_size[3]), .O(n23862) );
  ND2S U15036 ( .I1(n23932), .I2(n23900), .O(n23858) );
  ND2S U15037 ( .I1(n20606), .I2(n20524), .O(n16166) );
  OA22S U15038 ( .A1(n21254), .A2(n29503), .B1(n21467), .B2(n21259), .O(n20654) );
  ND2S U15039 ( .I1(n16963), .I2(n16962), .O(n16964) );
  NR2 U15040 ( .I1(n24692), .I2(n24614), .O(n24665) );
  NR2 U15041 ( .I1(n24681), .I2(n24692), .O(n24753) );
  ND2 U15042 ( .I1(n23974), .I2(n23961), .O(n24721) );
  ND2S U15043 ( .I1(n24748), .I2(n24105), .O(n24129) );
  NR2 U15044 ( .I1(n24350), .I2(n24669), .O(n24319) );
  NR2 U15045 ( .I1(n24646), .I2(n24692), .O(n24713) );
  ND2P U15046 ( .I1(n24665), .I2(n24721), .O(n24725) );
  NR3H U15047 ( .I1(n24099), .I2(n24098), .I3(n24097), .O(n24543) );
  NR2P U15048 ( .I1(n24099), .I2(n24111), .O(n24304) );
  NR3H U15049 ( .I1(n24013), .I2(n24098), .I3(n24097), .O(n24476) );
  ND2S U15050 ( .I1(n24517), .I2(n24516), .O(n29099) );
  ND2S U15051 ( .I1(n24542), .I2(n24515), .O(n24516) );
  ND2S U15052 ( .I1(n24517), .I2(n24196), .O(n29252) );
  ND2S U15053 ( .I1(n24622), .I2(n24515), .O(n24196) );
  ND2S U15054 ( .I1(n24517), .I2(n23987), .O(n28649) );
  ND2S U15055 ( .I1(n24670), .I2(n24515), .O(n23987) );
  AO12S U15056 ( .B1(n24476), .B2(n24670), .A1(n24510), .O(n28609) );
  AO12S U15057 ( .B1(n24476), .B2(n24585), .A1(n24510), .O(n29051) );
  AO12S U15058 ( .B1(n24543), .B2(n24542), .A1(n24541), .O(n29127) );
  AO12S U15059 ( .B1(n24543), .B2(n24585), .A1(n24541), .O(n29119) );
  AO12S U15060 ( .B1(n24543), .B2(n24346), .A1(n24541), .O(n29198) );
  ND2S U15061 ( .I1(n24517), .I2(n24406), .O(n28868) );
  ND2S U15062 ( .I1(n24515), .I2(n24727), .O(n24406) );
  AO12S U15063 ( .B1(n24476), .B2(n24542), .A1(n24510), .O(n29058) );
  AO12S U15064 ( .B1(n24277), .B2(n24444), .A1(n24541), .O(n28945) );
  AO12S U15065 ( .B1(n24476), .B2(n24346), .A1(n24510), .O(n29245) );
  AO12 U15066 ( .B1(n24463), .B2(n24585), .A1(n24462), .O(n29037) );
  ND2S U15067 ( .I1(n24298), .I2(n24517), .O(n28955) );
  ND2S U15068 ( .I1(n24304), .I2(n24622), .O(n24298) );
  AO12 U15069 ( .B1(n24134), .B2(n24515), .A1(n24462), .O(n28656) );
  AO12S U15070 ( .B1(n24543), .B2(n24444), .A1(n24541), .O(n28987) );
  AO12S U15071 ( .B1(n24543), .B2(n24727), .A1(n24541), .O(n28983) );
  ND2S U15072 ( .I1(n24244), .I2(n24517), .O(n28896) );
  ND2S U15073 ( .I1(n24250), .I2(n24622), .O(n24244) );
  AO12S U15074 ( .B1(n24476), .B2(n24727), .A1(n24510), .O(n28828) );
  ND2S U15075 ( .I1(n24517), .I2(n24200), .O(n29261) );
  ND2S U15076 ( .I1(n24346), .I2(n24515), .O(n24200) );
  AO12S U15077 ( .B1(n24304), .B2(n24444), .A1(n24541), .O(n28973) );
  AO12S U15078 ( .B1(n24476), .B2(n24444), .A1(n24541), .O(n28832) );
  ND2S U15079 ( .I1(n23859), .I2(n24332), .O(n13949) );
  HA1S U15080 ( .A(n21527), .B(n21526), .C(n21545), .S(n21528) );
  MUX2S U15081 ( .A(n29925), .B(n29924), .S(n29934), .O(n29955) );
  MUX2S U15082 ( .A(n29927), .B(n29926), .S(n29934), .O(n29953) );
  MUX2S U15083 ( .A(n29929), .B(n29928), .S(n29934), .O(n29951) );
  MUX2S U15084 ( .A(n29931), .B(n29930), .S(n29934), .O(n29949) );
  MUX2S U15085 ( .A(n29933), .B(n29932), .S(n29934), .O(n29947) );
  MUX2S U15086 ( .A(n29936), .B(n29935), .S(n29934), .O(n29945) );
  ND2S U15087 ( .I1(n13820), .I2(img[1224]), .O(n28286) );
  ND2S U15088 ( .I1(n13903), .I2(img[1226]), .O(n25434) );
  ND2S U15089 ( .I1(n13905), .I2(img[1239]), .O(n24460) );
  OR2S U15090 ( .I1(n21225), .I2(n20891), .O(n20859) );
  OR2S U15091 ( .I1(n13887), .I2(n29470), .O(n20858) );
  OA22S U15092 ( .A1(n21811), .A2(n21403), .B1(n21407), .B2(n21808), .O(n17961) );
  ND2S U15093 ( .I1(n20503), .I2(n22162), .O(n17695) );
  OR2S U15094 ( .I1(n21610), .I2(n28528), .O(n20726) );
  OR2S U15095 ( .I1(n29441), .I2(n27262), .O(n20725) );
  OA22S U15096 ( .A1(n22322), .A2(n21000), .B1(n20776), .B2(n23184), .O(n20698) );
  MOAI1S U15097 ( .A1(n15113), .A2(n30792), .B1(n15786), .B2(img[285]), .O(
        n15091) );
  MOAI1S U15098 ( .A1(n13894), .A2(n31005), .B1(n15786), .B2(img[293]), .O(
        n15115) );
  MOAI1S U15099 ( .A1(n15765), .A2(n30810), .B1(n13797), .B2(img[677]), .O(
        n15119) );
  OR2S U15100 ( .I1(n20903), .I2(n21411), .O(n20905) );
  AN2S U15101 ( .I1(n19059), .I2(n20780), .O(n20781) );
  OR2S U15102 ( .I1(n20892), .I2(n23185), .O(n20847) );
  MOAI1S U15103 ( .A1(n13850), .A2(n31896), .B1(n15809), .B2(img[1812]), .O(
        n15260) );
  MAO222S U15104 ( .A1(n21080), .B1(n28531), .C1(n28533), .O(n21084) );
  ND2S U15105 ( .I1(n21076), .I2(n21398), .O(n21015) );
  AN2S U15106 ( .I1(n21416), .I2(n29513), .O(n21271) );
  MOAI1S U15107 ( .A1(n13894), .A2(n30426), .B1(n15786), .B2(img[286]), .O(
        n15526) );
  MOAI1S U15108 ( .A1(n15113), .A2(n30300), .B1(n15786), .B2(img[318]), .O(
        n15550) );
  MOAI1S U15109 ( .A1(n15698), .A2(n30388), .B1(n17779), .B2(img[1878]), .O(
        n15456) );
  MOAI1S U15110 ( .A1(n13894), .A2(n31431), .B1(n15786), .B2(img[307]), .O(
        n14748) );
  MOAI1S U15111 ( .A1(n13894), .A2(n31408), .B1(n15786), .B2(img[267]), .O(
        n14723) );
  MOAI1S U15112 ( .A1(n13894), .A2(n31327), .B1(n15786), .B2(img[299]), .O(
        n14773) );
  ND2S U15113 ( .I1(n24768), .I2(n21416), .O(n21168) );
  AN2S U15114 ( .I1(n23839), .I2(n23846), .O(n21326) );
  OA22S U15115 ( .A1(n29441), .A2(n20892), .B1(n20899), .B2(n20740), .O(n20741) );
  AN2S U15116 ( .I1(n20137), .I2(n20136), .O(n13936) );
  ND2S U15117 ( .I1(n20161), .I2(n20363), .O(n20136) );
  ND3S U15118 ( .I1(n15287), .I2(n15286), .I3(n15285), .O(n15288) );
  ND2S U15119 ( .I1(n19059), .I2(n21412), .O(n21413) );
  OA22S U15120 ( .A1(n21259), .A2(n20788), .B1(n21254), .B2(n20784), .O(n20689) );
  INV1S U15121 ( .I(n21435), .O(n20797) );
  ND2S U15122 ( .I1(n20293), .I2(n19818), .O(n20296) );
  ND2S U15123 ( .I1(n20366), .I2(n20293), .O(n20295) );
  ND2S U15124 ( .I1(n19981), .I2(n19980), .O(n19982) );
  AN2S U15125 ( .I1(n19987), .I2(n20366), .O(n13944) );
  MOAI1S U15126 ( .A1(n13894), .A2(n30120), .B1(n15786), .B2(img[287]), .O(
        n15761) );
  MOAI1S U15127 ( .A1(n13894), .A2(n30182), .B1(n15786), .B2(img[319]), .O(
        n15788) );
  MOAI1S U15128 ( .A1(n15668), .A2(n30548), .B1(n15751), .B2(img[1842]), .O(
        n14315) );
  MOAI1S U15129 ( .A1(n14896), .A2(n30756), .B1(n15786), .B2(img[282]), .O(
        n14288) );
  MOAI1S U15130 ( .A1(n18141), .A2(n31180), .B1(n15751), .B2(img[1833]), .O(
        n14188) );
  MOAI1S U15131 ( .A1(n13894), .A2(n31115), .B1(n15786), .B2(img[281]), .O(
        n14121) );
  MOAI1S U15132 ( .A1(n13850), .A2(n31208), .B1(n15080), .B2(img[1993]), .O(
        n14110) );
  MOAI1S U15133 ( .A1(n15113), .A2(n31254), .B1(n15786), .B2(img[273]), .O(
        n14202) );
  MOAI1S U15134 ( .A1(n13894), .A2(n31655), .B1(n15786), .B2(img[264]), .O(
        n14656) );
  MOAI1S U15135 ( .A1(n13894), .A2(n31737), .B1(n15786), .B2(img[280]), .O(
        n14554) );
  MOAI1S U15136 ( .A1(n13894), .A2(n31722), .B1(n15786), .B2(img[304]), .O(
        n14605) );
  MOAI1S U15137 ( .A1(n17398), .A2(n17397), .B1(n17396), .B2(n19483), .O(
        n17402) );
  MOAI1S U15138 ( .A1(n17400), .A2(n17658), .B1(n17399), .B2(n20187), .O(
        n17401) );
  ND2P U15139 ( .I1(n21357), .I2(n21356), .O(n21377) );
  OR2S U15140 ( .I1(n21467), .I2(n23839), .O(n19440) );
  AN2S U15141 ( .I1(n23839), .I2(n21467), .O(n19439) );
  NR2P U15142 ( .I1(act_ptr[2]), .I2(act_ptr[1]), .O(n13988) );
  ND2S U15143 ( .I1(n20287), .I2(n20252), .O(n20253) );
  AN2S U15144 ( .I1(n19768), .I2(n19767), .O(n13906) );
  ND2S U15145 ( .I1(n19766), .I2(n20363), .O(n19767) );
  INV1 U15146 ( .I(n13766), .O(n20620) );
  MOAI1S U15147 ( .A1(n16228), .A2(n17397), .B1(n16238), .B2(n13843), .O(
        n15826) );
  OR2S U15148 ( .I1(i_col[3]), .I2(i_col[2]), .O(n14075) );
  ND2S U15149 ( .I1(n28547), .I2(A67_shift[252]), .O(n28548) );
  ND3S U15150 ( .I1(n26650), .I2(n26649), .I3(n26648), .O(n26662) );
  OR2S U15151 ( .I1(n26647), .I2(n28544), .O(n26648) );
  ND3S U15152 ( .I1(n25404), .I2(n28555), .I3(n25403), .O(n25407) );
  ND2S U15153 ( .I1(n28554), .I2(A67_shift[106]), .O(n25409) );
  ND2S U15154 ( .I1(n28547), .I2(A67_shift[232]), .O(n27900) );
  AN2S U15155 ( .I1(n28555), .I2(n27902), .O(n27903) );
  AO22S U15156 ( .A1(n28552), .A2(A67_shift[139]), .B1(n28553), .B2(
        A67_shift[11]), .O(n27270) );
  ND3S U15157 ( .I1(n27268), .I2(n28555), .I3(n27267), .O(n27269) );
  ND2S U15158 ( .I1(n28547), .I2(A67_shift[235]), .O(n27272) );
  AO22S U15159 ( .A1(n28552), .A2(A67_shift[155]), .B1(n28551), .B2(
        A67_shift[219]), .O(n27277) );
  ND3S U15160 ( .I1(n27275), .I2(n27274), .I3(n28540), .O(n27276) );
  ND2S U15161 ( .I1(n20608), .I2(n19818), .O(n16201) );
  ND3S U15162 ( .I1(n16206), .I2(n16205), .I3(n16204), .O(n16210) );
  BUF2 U15163 ( .I(n16200), .O(n22923) );
  INV2 U15164 ( .I(n16188), .O(n19661) );
  ND2S U15165 ( .I1(n20809), .I2(n24701), .O(n13999) );
  ND2 U15166 ( .I1(n23665), .I2(n13939), .O(n23797) );
  ND2S U15167 ( .I1(n24722), .I2(n24664), .O(n24735) );
  NR2 U15168 ( .I1(n24692), .I2(n24476), .O(n24479) );
  OR2S U15169 ( .I1(n24705), .I2(n24707), .O(n24764) );
  AN2S U15170 ( .I1(n24707), .I2(n24706), .O(n24763) );
  NR2 U15171 ( .I1(n24692), .I2(n24304), .O(n24293) );
  NR2P U15172 ( .I1(n24692), .I2(n23909), .O(n24957) );
  NR2 U15173 ( .I1(n24697), .I2(n24097), .O(n23909) );
  NR2P U15174 ( .I1(n24692), .I2(n23968), .O(n24732) );
  INV1S U15175 ( .I(n24659), .O(n23968) );
  NR2 U15176 ( .I1(n24673), .I2(n24692), .O(n24744) );
  INV1S U15177 ( .I(n24668), .O(n24740) );
  ND2S U15178 ( .I1(addr[7]), .I2(addr[6]), .O(n13950) );
  NR2 U15179 ( .I1(n24563), .I2(n24957), .O(n29136) );
  AO12S U15180 ( .B1(n24665), .B2(n24509), .A1(n24682), .O(n28645) );
  AO12S U15181 ( .B1(n24665), .B2(n24664), .A1(n24682), .O(n29318) );
  NR2 U15182 ( .I1(n24682), .I2(n24038), .O(n28686) );
  NR2 U15183 ( .I1(n24682), .I2(n24084), .O(n28743) );
  NR2 U15184 ( .I1(n24682), .I2(n23939), .O(n28605) );
  NR2 U15185 ( .I1(n24682), .I2(n24653), .O(n29306) );
  ND2S U15186 ( .I1(n24501), .I2(n24495), .O(n29081) );
  ND2S U15187 ( .I1(n24500), .I2(n24735), .O(n24501) );
  NR2 U15188 ( .I1(n24159), .I2(n24319), .O(n29214) );
  NR2 U15189 ( .I1(n24175), .I2(n24319), .O(n29221) );
  NR2 U15190 ( .I1(n24217), .I2(n24319), .O(n29201) );
  NR2 U15191 ( .I1(n24140), .I2(n24319), .O(n29283) );
  NR2 U15192 ( .I1(n24529), .I2(n24957), .O(n29030) );
  NR2 U15193 ( .I1(n24006), .I2(n24957), .O(n28587) );
  NR2 U15194 ( .I1(n24184), .I2(n24957), .O(n29276) );
  ND2S U15195 ( .I1(n24744), .I2(n24694), .O(n24625) );
  ND2S U15196 ( .I1(n24479), .I2(n24758), .O(n24469) );
  OA12S U15197 ( .B1(n24238), .B2(n24105), .A1(n24748), .O(n28693) );
  OA12S U15198 ( .B1(n24238), .B2(n24023), .A1(n24495), .O(n28679) );
  NR2 U15199 ( .I1(n24229), .I2(n24335), .O(n29007) );
  NR2 U15200 ( .I1(n24229), .I2(n24238), .O(n28906) );
  NR2 U15201 ( .I1(n24229), .I2(n24744), .O(n29423) );
  NR2 U15202 ( .I1(n24229), .I2(n24753), .O(n29430) );
  NR2 U15203 ( .I1(n24229), .I2(n24732), .O(n29409) );
  NR2 U15204 ( .I1(n24319), .I2(n24251), .O(n28899) );
  ND2S U15205 ( .I1(n24736), .I2(n24689), .O(n29383) );
  OA12S U15206 ( .B1(n24266), .B2(n24023), .A1(n24495), .O(n28708) );
  NR2 U15207 ( .I1(n23916), .I2(n24682), .O(n28590) );
  NR2 U15208 ( .I1(n24641), .I2(n24682), .O(n29289) );
  NR2 U15209 ( .I1(n24440), .I2(n24379), .O(n28835) );
  NR2 U15210 ( .I1(n24409), .I2(n24440), .O(n28875) );
  NR2 U15211 ( .I1(n24229), .I2(n24479), .O(n28824) );
  NR2 U15212 ( .I1(n24425), .I2(n24957), .O(n28807) );
  NR2 U15213 ( .I1(n24647), .I2(n24682), .O(n29300) );
  NR2 U15214 ( .I1(n24674), .I2(n24682), .O(n29324) );
  NR2 U15215 ( .I1(n24683), .I2(n24682), .O(n29331) );
  NR2 U15216 ( .I1(n24578), .I2(n24957), .O(n29139) );
  ND2S U15217 ( .I1(n24546), .I2(n24694), .O(n24308) );
  AO12S U15218 ( .B1(n24250), .B2(n24585), .A1(n24510), .O(n28676) );
  AO12S U15219 ( .B1(n24277), .B2(n24585), .A1(n24510), .O(n28705) );
  ND2S U15220 ( .I1(n24293), .I2(n24748), .O(n24091) );
  OA12S U15221 ( .B1(n24546), .B2(n24023), .A1(n24495), .O(n29122) );
  ND2S U15222 ( .I1(n24449), .I2(n24495), .O(n29021) );
  ND2S U15223 ( .I1(n24500), .I2(n24689), .O(n24449) );
  OA12S U15224 ( .B1(n24490), .B2(n24726), .A1(n24725), .O(n29067) );
  NR2 U15225 ( .I1(n24319), .I2(n24318), .O(n29192) );
  NR2 U15226 ( .I1(n24636), .I2(n24957), .O(n29339) );
  NR2 U15227 ( .I1(n24958), .I2(n24957), .O(n29536) );
  NR2 U15228 ( .I1(n24105), .I2(n24957), .O(n28584) );
  ND2S U15229 ( .I1(n24293), .I2(n24694), .O(n24294) );
  OA12S U15230 ( .B1(n24546), .B2(n24105), .A1(n24748), .O(n28764) );
  AO12S U15231 ( .B1(n24351), .B2(n24585), .A1(n24510), .O(n28775) );
  NR2 U15232 ( .I1(n24229), .I2(n24266), .O(n28936) );
  NR2 U15233 ( .I1(n24229), .I2(n24293), .O(n28965) );
  OAI12HS U15234 ( .B1(n24105), .B2(n24520), .A1(n24748), .O(n28652) );
  NR2 U15235 ( .I1(n24319), .I2(n24305), .O(n28958) );
  NR2 U15236 ( .I1(n24440), .I2(n24254), .O(n28948) );
  NR2 U15237 ( .I1(n24440), .I2(n24280), .O(n28976) );
  NR2 U15238 ( .I1(n24229), .I2(n24546), .O(n28979) );
  NR2 U15239 ( .I1(n24440), .I2(n24439), .O(n28990) );
  NR2 U15240 ( .I1(n24612), .I2(n24957), .O(n29342) );
  NR2 U15241 ( .I1(n24229), .I2(n24713), .O(n29395) );
  AO12S U15242 ( .B1(n24543), .B2(n24622), .A1(n24541), .O(n29189) );
  ND2S U15243 ( .I1(n24271), .I2(n24517), .O(n28926) );
  ND2S U15244 ( .I1(n24277), .I2(n24622), .O(n24271) );
  AO12S U15245 ( .B1(n24476), .B2(n24622), .A1(n24510), .O(n29237) );
  ND2S U15246 ( .I1(n24351), .I2(n24727), .O(n24331) );
  AO12S U15247 ( .B1(n24543), .B2(n24766), .A1(n24726), .O(n28757) );
  ND2S U15248 ( .I1(n24758), .I2(n24744), .O(n24575) );
  ND3S U15249 ( .I1(n28569), .I2(n28568), .I3(n28567), .O(n28570) );
  AOI12HP U15250 ( .B1(n26670), .B2(n28575), .A1(n26669), .O(n27170) );
  ND3S U15251 ( .I1(n26666), .I2(n26665), .I3(n26664), .O(n26667) );
  ND2S U15252 ( .I1(n24790), .I2(n24789), .O(n24791) );
  ND3S U15253 ( .I1(n23888), .I2(n23887), .I3(n23886), .O(n23889) );
  AO12 U15254 ( .B1(n24351), .B2(n24444), .A1(n24541), .O(n29015) );
  ND2S U15255 ( .I1(n25416), .I2(n25415), .O(n25417) );
  ND3S U15256 ( .I1(n27285), .I2(n27284), .I3(n27283), .O(n27286) );
  AO12S U15257 ( .B1(n24304), .B2(n24585), .A1(n24510), .O(n28733) );
  ND3S U15258 ( .I1(n26035), .I2(n26034), .I3(n26033), .O(n26036) );
  AO12 U15259 ( .B1(n24515), .B2(n24444), .A1(n24541), .O(n28872) );
  ND2S U15260 ( .I1(n24341), .I2(n24517), .O(n28997) );
  ND2S U15261 ( .I1(n24351), .I2(n24622), .O(n24341) );
  AO12 U15262 ( .B1(n24351), .B2(n24542), .A1(n24263), .O(n28782) );
  AO12 U15263 ( .B1(n24277), .B2(n24134), .A1(n24462), .O(n28726) );
  NR2 U15264 ( .I1(n24511), .I2(n24510), .O(n29091) );
  AO12S U15265 ( .B1(n24543), .B2(n24134), .A1(n24541), .O(n28768) );
  AO12S U15266 ( .B1(n24250), .B2(n24444), .A1(n24541), .O(n28916) );
  ND2S U15267 ( .I1(n29521), .I2(n21602), .O(n21603) );
  ND2S U15268 ( .I1(n23038), .I2(n23037), .O(n23132) );
  ND2S U15269 ( .I1(n23326), .I2(n23325), .O(n23385) );
  ND2S U15270 ( .I1(n22516), .I2(n22515), .O(n22614) );
  ND2S U15271 ( .I1(n22512), .I2(n22511), .O(n22625) );
  ND2S U15272 ( .I1(n21964), .I2(n21963), .O(n21999) );
  ND2S U15273 ( .I1(n22216), .I2(n22215), .O(n22251) );
  ND2S U15274 ( .I1(c_s[0]), .I2(n14029), .O(n14012) );
  MAO222 U15275 ( .A1(n29923), .B1(rgb_value[15]), .C1(n29922), .O(n29934) );
  MAO222 U15276 ( .A1(n29925), .B1(rgb_value[14]), .C1(n29921), .O(n29922) );
  MAO222 U15277 ( .A1(n29927), .B1(rgb_value[13]), .C1(n29920), .O(n29921) );
  MAO222 U15278 ( .A1(rgb_value[7]), .B1(n29943), .C1(n29942), .O(n29956) );
  MAO222 U15279 ( .A1(n29955), .B1(rgb_value[6]), .C1(n29941), .O(n29942) );
  MAO222 U15280 ( .A1(rgb_value[5]), .B1(n29953), .C1(n29940), .O(n29941) );
  MAO222 U15281 ( .A1(n29951), .B1(rgb_value[4]), .C1(n29939), .O(n29940) );
  ND2S U15282 ( .I1(n13770), .I2(img[1482]), .O(n25472) );
  ND2S U15283 ( .I1(n13905), .I2(img[1489]), .O(n26977) );
  ND2S U15284 ( .I1(n13905), .I2(img[1507]), .O(n27807) );
  ND2S U15285 ( .I1(n29124), .I2(img[1490]), .O(n25624) );
  ND2S U15286 ( .I1(n13820), .I2(img[1889]), .O(n26736) );
  ND2S U15287 ( .I1(n29124), .I2(img[1888]), .O(n27930) );
  ND2S U15288 ( .I1(n29124), .I2(img[1890]), .O(n25762) );
  ND2S U15289 ( .I1(n29124), .I2(img[1656]), .O(n28044) );
  ND2S U15290 ( .I1(n13905), .I2(img[1354]), .O(n25445) );
  ND2S U15291 ( .I1(n29124), .I2(img[1216]), .O(n27920) );
  ND2S U15292 ( .I1(n13900), .I2(img[1264]), .O(n28283) );
  ND2S U15293 ( .I1(n29258), .I2(img[1266]), .O(n25431) );
  ND2S U15294 ( .I1(n29124), .I2(img[1500]), .O(n29259) );
  ND2S U15295 ( .I1(n29124), .I2(img[1404]), .O(n28830) );
  ND2S U15296 ( .I1(n13820), .I2(img[1252]), .O(n29209) );
  ND2S U15297 ( .I1(n13904), .I2(img[1495]), .O(n24513) );
  ND2S U15298 ( .I1(n29124), .I2(img[1247]), .O(n24155) );
  ND2S U15299 ( .I1(n13903), .I2(img[1367]), .O(n24474) );
  ND2S U15300 ( .I1(n13820), .I2(img[1103]), .O(n24101) );
  ND2S U15301 ( .I1(n13819), .I2(img[1263]), .O(n24457) );
  ND2S U15302 ( .I1(n13820), .I2(img[1494]), .O(n25293) );
  ND2S U15303 ( .I1(n29124), .I2(img[1497]), .O(n26870) );
  ND2S U15304 ( .I1(n29124), .I2(img[1502]), .O(n25155) );
  ND2S U15305 ( .I1(n13820), .I2(img[1273]), .O(n26681) );
  ND2S U15306 ( .I1(n13819), .I2(img[1254]), .O(n25116) );
  ND2S U15307 ( .I1(n13901), .I2(img[1238]), .O(n25322) );
  ND2S U15308 ( .I1(n29124), .I2(img[1406]), .O(n24819) );
  ND2S U15309 ( .I1(n13903), .I2(img[1134]), .O(n25307) );
  ND2S U15310 ( .I1(n13820), .I2(img[1366]), .O(n25283) );
  ND2S U15311 ( .I1(n13820), .I2(img[1385]), .O(n26955) );
  ND2S U15312 ( .I1(n13820), .I2(img[1094]), .O(n24921) );
  ND2S U15313 ( .I1(n13820), .I2(img[1097]), .O(n27154) );
  ND2S U15314 ( .I1(n13820), .I2(img[1102]), .O(n25083) );
  ND2S U15315 ( .I1(n13820), .I2(img[1113]), .O(n26889) );
  ND2S U15316 ( .I1(n13770), .I2(img[1118]), .O(n25175) );
  ND2S U15317 ( .I1(n13820), .I2(img[1475]), .O(n27528) );
  ND2S U15318 ( .I1(n13820), .I2(img[1491]), .O(n27340) );
  ND2S U15319 ( .I1(n13820), .I2(img[1403]), .O(n27506) );
  ND2S U15320 ( .I1(n13820), .I2(img[1275]), .O(n27496) );
  ND2S U15321 ( .I1(n13820), .I2(img[1099]), .O(n27711) );
  ND2S U15322 ( .I1(n13820), .I2(img[1107]), .O(n27422) );
  ND2S U15323 ( .I1(n13819), .I2(img[1355]), .O(n27664) );
  ND2S U15324 ( .I1(n13820), .I2(img[1363]), .O(n27313) );
  ND2S U15325 ( .I1(n13820), .I2(img[1235]), .O(n27303) );
  ND2S U15326 ( .I1(n13820), .I2(img[1496]), .O(n28397) );
  ND2S U15327 ( .I1(n13905), .I2(img[1498]), .O(n25912) );
  ND2S U15328 ( .I1(n13820), .I2(img[1634]), .O(n25802) );
  ND2S U15329 ( .I1(n13900), .I2(img[1400]), .O(n27974) );
  ND2S U15330 ( .I1(n29124), .I2(img[1786]), .O(n25792) );
  ND2S U15331 ( .I1(n13820), .I2(img[1114]), .O(n25931) );
  ND2S U15332 ( .I1(n13820), .I2(img[1146]), .O(n25823) );
  ND2S U15333 ( .I1(n13905), .I2(img[1520]), .O(n28321) );
  ND2S U15334 ( .I1(n13819), .I2(img[1373]), .O(n26065) );
  ND2S U15335 ( .I1(n13820), .I2(img[1117]), .O(n26177) );
  ND2S U15336 ( .I1(n13905), .I2(img[1478]), .O(n24840) );
  ND2S U15337 ( .I1(n13903), .I2(img[1374]), .O(n25129) );
  ND2S U15338 ( .I1(n13819), .I2(img[1907]), .O(n27356) );
  ND2S U15339 ( .I1(n13902), .I2(img[1349]), .O(n26377) );
  OR2 U15340 ( .I1(n21545), .I2(n21536), .O(gray_avg[7]) );
  OR2 U15341 ( .I1(n21573), .I2(n21564), .O(gray_avg[5]) );
  OR2 U15342 ( .I1(n23440), .I2(n21593), .O(gray_avg[3]) );
  OR2S U15343 ( .I1(n23465), .I2(n23458), .O(gray_avg[1]) );
  HA1S U15344 ( .A(PE_mul[35]), .B(PE_mul[3]), .C(n29575), .S(n29568) );
  AO12S U15345 ( .B1(n29470), .B2(n29463), .A1(n20811), .O(n20814) );
  OR2S U15346 ( .I1(n22668), .I2(n29470), .O(n20813) );
  OR2S U15347 ( .I1(n23188), .I2(n21394), .O(n20994) );
  OR2S U15348 ( .I1(n21399), .I2(n21398), .O(n21401) );
  MOAI1S U15349 ( .A1(n15698), .A2(n30324), .B1(n13828), .B2(img[1830]), .O(
        n15467) );
  INV2 U15350 ( .I(i_row[1]), .O(n14043) );
  INV2 U15351 ( .I(n14112), .O(n16016) );
  BUF1S U15352 ( .I(n19710), .O(n18892) );
  BUF1S U15353 ( .I(n19710), .O(n19031) );
  BUF1S U15354 ( .I(n19710), .O(n19313) );
  MOAI1S U15355 ( .A1(n14896), .A2(n30959), .B1(n15786), .B2(img[309]), .O(
        n14991) );
  MOAI1S U15356 ( .A1(n15113), .A2(n30931), .B1(n15786), .B2(img[301]), .O(
        n14942) );
  MOAI1S U15357 ( .A1(n15780), .A2(n30909), .B1(n15809), .B2(img[1917]), .O(
        n14963) );
  MOAI1S U15358 ( .A1(n14896), .A2(n30851), .B1(n15786), .B2(img[277]), .O(
        n15041) );
  ND2S U15359 ( .I1(n29461), .I2(n29475), .O(n18668) );
  OR2S U15360 ( .I1(n21658), .I2(n29470), .O(n20737) );
  OA22S U15361 ( .A1(n20863), .A2(n20899), .B1(n20903), .B2(n21245), .O(n20864) );
  ND2P U15362 ( .I1(i_row[2]), .I2(i_row[3]), .O(n14033) );
  OR2S U15363 ( .I1(n21808), .I2(n20899), .O(n19617) );
  MOAI1S U15364 ( .A1(n15780), .A2(n31936), .B1(n17088), .B2(img[1380]), .O(
        n15283) );
  INV2 U15365 ( .I(n14266), .O(n16326) );
  OR2S U15366 ( .I1(n29489), .I2(n22667), .O(n21119) );
  OA22S U15367 ( .A1(n22920), .A2(n24768), .B1(n26012), .B2(n22922), .O(n21122) );
  OAI112HS U15368 ( .C1(n21403), .C2(n22932), .A1(n21251), .B1(n21250), .O(
        n21252) );
  OR2S U15369 ( .I1(n21407), .I2(n28527), .O(n21409) );
  ND2S U15370 ( .I1(n17962), .I2(n17961), .O(n17964) );
  OR2S U15371 ( .I1(n21392), .I2(n23845), .O(n20732) );
  BUF1 U15372 ( .I(n19710), .O(n19266) );
  BUF3 U15373 ( .I(n22928), .O(n20193) );
  BUF6 U15374 ( .I(n14077), .O(n18297) );
  INV3 U15375 ( .I(n18155), .O(n15277) );
  MOAI1S U15376 ( .A1(n16720), .A2(n13766), .B1(n16719), .B2(n17938), .O(
        n16724) );
  NR2P U15377 ( .I1(n14033), .I2(n14058), .O(n16003) );
  INV2 U15378 ( .I(n29448), .O(n21117) );
  MOAI1S U15379 ( .A1(n14896), .A2(n31491), .B1(n15786), .B2(img[283]), .O(
        n14847) );
  MAO222S U15380 ( .A1(n21158), .B1(n25391), .C1(n29497), .O(n21165) );
  ND2S U15381 ( .I1(n27262), .I2(n29455), .O(n21161) );
  AN2S U15382 ( .I1(n23845), .I2(n23839), .O(n21171) );
  ND2S U15383 ( .I1(n21416), .I2(n29503), .O(n19238) );
  OR2S U15384 ( .I1(n19461), .I2(n23839), .O(n20911) );
  AN2S U15385 ( .I1(n23839), .I2(n19461), .O(n20910) );
  AN2S U15386 ( .I1(n23839), .I2(n20788), .O(n20789) );
  OR2S U15387 ( .I1(n22671), .I2(n20892), .O(n20818) );
  AN2S U15388 ( .I1(n22412), .I2(n21340), .O(n20836) );
  INV2 U15389 ( .I(n21479), .O(n21474) );
  BUF3 U15390 ( .I(n19642), .O(n17376) );
  OR2S U15391 ( .I1(n21660), .I2(n21595), .O(n20398) );
  AO12S U15392 ( .B1(n20535), .B2(n28528), .A1(n20378), .O(n13937) );
  MOAI1S U15393 ( .A1(n17940), .A2(n13927), .B1(n17936), .B2(n21062), .O(
        n15367) );
  MOAI1S U15394 ( .A1(n15363), .A2(n19462), .B1(n17929), .B2(n17875), .O(
        n15365) );
  MOAI1S U15395 ( .A1(n17930), .A2(n13945), .B1(n17932), .B2(n20263), .O(
        n15364) );
  AN2S U15396 ( .I1(n23839), .I2(n20855), .O(n21277) );
  ND3S U15397 ( .I1(n20284), .I2(n20283), .I3(n20282), .O(n20285) );
  ND2S U15398 ( .I1(n20366), .I2(n20281), .O(n20283) );
  AO22S U15399 ( .A1(n20063), .A2(n20685), .B1(n19818), .B2(n19987), .O(n13924) );
  ND2S U15400 ( .I1(n19696), .I2(n20363), .O(n19697) );
  BUF1S U15401 ( .I(n19710), .O(n19253) );
  MOAI1S U15402 ( .A1(n16491), .A2(n17397), .B1(n16493), .B2(n17938), .O(
        n15590) );
  MOAI1S U15403 ( .A1(n16488), .A2(n13947), .B1(n16476), .B2(n20629), .O(
        n15589) );
  OA22S U15404 ( .A1(n15142), .A2(n17421), .B1(n17412), .B2(n19462), .O(n14493) );
  MOAI1S U15405 ( .A1(n17400), .A2(n16468), .B1(n17403), .B2(n17931), .O(
        n14496) );
  MOAI1S U15406 ( .A1(n14896), .A2(n30728), .B1(n15786), .B2(img[290]), .O(
        n14338) );
  ND3S U15407 ( .I1(n14302), .I2(n14301), .I3(n14300), .O(n14306) );
  MOAI1S U15408 ( .A1(n15631), .A2(n30658), .B1(n19642), .B2(img[250]), .O(
        n14404) );
  INV2 U15409 ( .I(n19642), .O(n14092) );
  MOAI1S U15410 ( .A1(n17930), .A2(n13766), .B1(n17929), .B2(n17928), .O(
        n17935) );
  MOAI1S U15411 ( .A1(n17916), .A2(n13946), .B1(n17915), .B2(n13830), .O(
        n17927) );
  MOAI1S U15412 ( .A1(n17412), .A2(n13844), .B1(n17411), .B2(n13847), .O(
        n17416) );
  ND2S U15413 ( .I1(n17947), .I2(n17946), .O(n17948) );
  INV2 U15414 ( .I(n20385), .O(n20685) );
  ND2S U15415 ( .I1(img_size[1]), .I2(n23900), .O(n23860) );
  ND3S U15416 ( .I1(n19936), .I2(n19935), .I3(n19934), .O(n20012) );
  HA1S U15417 ( .A(n29555), .B(n29554), .C(n29557), .S(n29559) );
  OR2S U15418 ( .I1(n20788), .I2(n22410), .O(n20747) );
  ND2S U15419 ( .I1(n20259), .I2(n22923), .O(n16258) );
  ND2S U15420 ( .I1(n20259), .I2(n19818), .O(n16256) );
  ND3S U15421 ( .I1(n20274), .I2(n20273), .I3(n20272), .O(n20275) );
  ND3S U15422 ( .I1(n20266), .I2(n20265), .I3(n20264), .O(n20276) );
  ND2S U15423 ( .I1(n22055), .I2(n21340), .O(n21341) );
  ND2S U15424 ( .I1(n23839), .I2(n21449), .O(n21420) );
  MOAI1S U15425 ( .A1(n16241), .A2(n13946), .B1(n16227), .B2(n20439), .O(
        n15820) );
  MOAI1S U15426 ( .A1(n17659), .A2(n16468), .B1(n17669), .B2(n20263), .O(
        n14931) );
  MOAI1S U15427 ( .A1(n17657), .A2(n13946), .B1(n17663), .B2(n17938), .O(
        n14930) );
  MOAI1S U15428 ( .A1(n17670), .A2(n13947), .B1(n17677), .B2(n20406), .O(
        n14935) );
  MOAI1S U15429 ( .A1(n17675), .A2(n17656), .B1(n17671), .B2(n21062), .O(
        n14933) );
  MOAI1S U15430 ( .A1(n14076), .A2(n19462), .B1(n16947), .B2(n13846), .O(
        n14104) );
  NR2 U15431 ( .I1(n15665), .I2(n15664), .O(n16228) );
  ND3S U15432 ( .I1(n14291), .I2(n14290), .I3(n14289), .O(n14298) );
  MOAI1S U15433 ( .A1(n16933), .A2(n19462), .B1(n16932), .B2(n17938), .O(
        n16937) );
  MOAI1S U15434 ( .A1(n17159), .A2(n15142), .B1(n17158), .B2(n21062), .O(
        n17163) );
  MOAI1S U15435 ( .A1(n17172), .A2(n17397), .B1(n17171), .B2(n13830), .O(
        n17176) );
  MOAI1S U15436 ( .A1(n17174), .A2(n17658), .B1(n17173), .B2(n17938), .O(
        n17175) );
  OR2S U15437 ( .I1(n19554), .I2(n19574), .O(n19555) );
  NR2T U15438 ( .I1(n13844), .I2(n18133), .O(n19818) );
  INV1S U15439 ( .I(n23870), .O(n23740) );
  ND2S U15440 ( .I1(n13986), .I2(act[3]), .O(n13971) );
  FA1S U15441 ( .A(rgb_value[5]), .B(rgb_value[21]), .CI(rgb_value[13]), .CO(
        n21519), .S(n21518) );
  FA1S U15442 ( .A(rgb_value[4]), .B(rgb_value[20]), .CI(rgb_value[12]), .CO(
        n21517), .S(n21514) );
  FA1S U15443 ( .A(rgb_value[3]), .B(rgb_value[19]), .CI(rgb_value[11]), .CO(
        n21513), .S(n21512) );
  FA1S U15444 ( .A(rgb_value[2]), .B(rgb_value[18]), .CI(rgb_value[10]), .CO(
        n21511), .S(n21510) );
  ND2S U15445 ( .I1(n23908), .I2(n23974), .O(n24697) );
  ND2S U15446 ( .I1(col[2]), .I2(col[3]), .O(n24139) );
  AO22S U15447 ( .A1(n28552), .A2(A67_shift[159]), .B1(n28553), .B2(
        A67_shift[31]), .O(n23877) );
  ND2S U15448 ( .I1(n28547), .I2(A67_shift[255]), .O(n23879) );
  AO22S U15449 ( .A1(n28552), .A2(A67_shift[143]), .B1(n28551), .B2(
        A67_shift[207]), .O(n23866) );
  ND3S U15450 ( .I1(n23864), .I2(n28555), .I3(n23863), .O(n23865) );
  AO22S U15451 ( .A1(n28552), .A2(A67_shift[157]), .B1(n28553), .B2(
        A67_shift[29]), .O(n26027) );
  ND3S U15452 ( .I1(n26025), .I2(n26024), .I3(n28540), .O(n26026) );
  ND2S U15453 ( .I1(n28547), .I2(A67_shift[253]), .O(n26029) );
  AO22S U15454 ( .A1(n28552), .A2(A67_shift[141]), .B1(n28553), .B2(
        A67_shift[13]), .O(n26020) );
  OR2S U15455 ( .I1(n24032), .I2(n24700), .O(n24042) );
  NR2 U15456 ( .I1(n24097), .I2(n24112), .O(n23982) );
  INV2 U15457 ( .I(n24012), .O(n24097) );
  NR2 U15458 ( .I1(n24097), .I2(n24051), .O(n23961) );
  MOAI1S U15459 ( .A1(n17672), .A2(n20421), .B1(n17671), .B2(n13846), .O(
        n17673) );
  MOAI1S U15460 ( .A1(n17670), .A2(n13946), .B1(n17669), .B2(n20406), .O(
        n17674) );
  ND2S U15461 ( .I1(n19939), .I2(n19818), .O(n16438) );
  ND3S U15462 ( .I1(n20572), .I2(n20571), .I3(n13822), .O(n20576) );
  MOAI1S U15463 ( .A1(n20587), .A2(n20586), .B1(n20585), .B2(n20263), .O(
        n20591) );
  ND2S U15464 ( .I1(n20563), .I2(n20562), .O(n20564) );
  ND2S U15465 ( .I1(n19924), .I2(n19923), .O(n19925) );
  HA1S U15466 ( .A(n29557), .B(n29556), .C(n29874), .S(n29810) );
  OAI12HS U15467 ( .B1(n13968), .B2(n13967), .A1(n13966), .O(n23852) );
  ND2S U15468 ( .I1(n19452), .I2(n18142), .O(n22916) );
  INV2 U15469 ( .I(n21085), .O(n23848) );
  ND2S U15470 ( .I1(n19602), .I2(n18142), .O(n22938) );
  OA22S U15471 ( .A1(n21669), .A2(n21449), .B1(n17965), .B2(n21653), .O(n20762) );
  OA22S U15472 ( .A1(n22661), .A2(n21449), .B1(n22171), .B2(n21191), .O(n21192) );
  MAO222S U15473 ( .A1(n21435), .B1(n21438), .C1(n21436), .O(n21433) );
  AN2 U15474 ( .I1(n19603), .I2(n16464), .O(n20252) );
  INV3 U15475 ( .I(n13844), .O(n20969) );
  BUF4 U15476 ( .I(n15579), .O(n21254) );
  OR2S U15477 ( .I1(n19575), .I2(n19574), .O(n19576) );
  NR2T U15478 ( .I1(n18141), .I2(n19700), .O(n19608) );
  INV4 U15479 ( .I(n19661), .O(n20364) );
  HA1S U15480 ( .A(rgb_value[1]), .B(rgb_value[17]), .C(n21509), .S(n21507) );
  ND3S U15481 ( .I1(n24012), .I2(n23967), .I3(n23974), .O(n24659) );
  AN2S U15482 ( .I1(n24015), .I2(n24014), .O(n24568) );
  ND3S U15483 ( .I1(n28539), .I2(n28538), .I3(n28537), .O(n28563) );
  ND3S U15484 ( .I1(n28559), .I2(n28558), .I3(n28557), .O(n28560) );
  ND2S U15485 ( .I1(n28549), .I2(n28548), .O(n28561) );
  ND2S U15486 ( .I1(n26644), .I2(n26643), .O(n26663) );
  ND3S U15487 ( .I1(n26659), .I2(n26658), .I3(n26657), .O(n26660) );
  ND3S U15488 ( .I1(n24778), .I2(n24777), .I3(n24776), .O(n24787) );
  ND2S U15489 ( .I1(n23882), .I2(n23881), .O(n23890) );
  ND3S U15490 ( .I1(n23873), .I2(n23872), .I3(n23871), .O(n23882) );
  ND3S U15491 ( .I1(n23880), .I2(n23879), .I3(n23878), .O(n23881) );
  ND2S U15492 ( .I1(n28547), .I2(A67_shift[239]), .O(n23872) );
  ND3S U15493 ( .I1(n25411), .I2(n25410), .I3(n25409), .O(n25412) );
  ND3S U15494 ( .I1(n27896), .I2(n27895), .I3(n27894), .O(n27909) );
  ND3S U15495 ( .I1(n27905), .I2(n27904), .I3(n27903), .O(n27906) );
  ND2S U15496 ( .I1(n27901), .I2(n27900), .O(n27907) );
  ND2S U15497 ( .I1(n27282), .I2(n27281), .O(n27287) );
  ND3S U15498 ( .I1(n27273), .I2(n27272), .I3(n27271), .O(n27282) );
  ND2S U15499 ( .I1(n28547), .I2(A67_shift[251]), .O(n27279) );
  ND2S U15500 ( .I1(n26032), .I2(n26031), .O(n26037) );
  ND3S U15501 ( .I1(n26023), .I2(n26022), .I3(n26021), .O(n26032) );
  ND3S U15502 ( .I1(n26030), .I2(n26029), .I3(n26028), .O(n26031) );
  ND2S U15503 ( .I1(n28547), .I2(A67_shift[237]), .O(n26022) );
  NR2 U15504 ( .I1(n23927), .I2(n24517), .O(n24510) );
  NR2 U15505 ( .I1(n23926), .I2(n24541), .O(n24517) );
  NR2 U15506 ( .I1(n24332), .I2(n24034), .O(n23926) );
  BUF2 U15507 ( .I(n19700), .O(n21654) );
  INV1 U15508 ( .I(n21079), .O(n29443) );
  ND2 U15509 ( .I1(n22921), .I2(n20809), .O(n19058) );
  INV1 U15510 ( .I(n21399), .O(n29491) );
  INV2 U15511 ( .I(n21076), .O(n29484) );
  AO12S U15512 ( .B1(n29842), .B2(n29841), .A1(n29777), .O(n29808) );
  HA1S U15513 ( .A(n29874), .B(n29873), .C(n29807), .S(n29908) );
  INV2 U15514 ( .I(i_row[0]), .O(n23824) );
  ND2 U15515 ( .I1(n16185), .I2(n16184), .O(n16186) );
  NR2 U15516 ( .I1(n16179), .I2(n23797), .O(n16185) );
  ND2S U15517 ( .I1(n14030), .I2(n23565), .O(n23572) );
  AOI12HS U15518 ( .B1(n16226), .B2(n20364), .A1(n16203), .O(n16213) );
  ND2S U15519 ( .I1(n16202), .I2(n16201), .O(n16203) );
  NR2 U15520 ( .I1(n22923), .I2(n13822), .O(n19438) );
  OAI22S U15521 ( .A1(n18489), .A2(n19235), .B1(n18489), .B2(n19661), .O(
        n18491) );
  HA1S U15522 ( .A(n22724), .B(n22723), .C(n22721), .S(n22733) );
  HA1S U15523 ( .A(n23240), .B(n23239), .C(n23237), .S(n23252) );
  HA1S U15524 ( .A(n23246), .B(n23245), .C(n23241), .S(n23250) );
  HA1S U15525 ( .A(n22477), .B(n22476), .C(n22472), .S(n22481) );
  HA1S U15526 ( .A(n21865), .B(n21864), .C(n21862), .S(n21874) );
  HA1S U15527 ( .A(n22114), .B(n22113), .C(n22111), .S(n22126) );
  ND2S U15528 ( .I1(n23718), .I2(n23717), .O(n23719) );
  INV1S U15529 ( .I(n30039), .O(n23730) );
  OA12S U15530 ( .B1(n14023), .B2(n14022), .A1(n31997), .O(n14024) );
  OR2S U15531 ( .I1(set_cnt[1]), .I2(set_cnt[2]), .O(n14022) );
  MAO222S U15532 ( .A1(n29929), .B1(rgb_value[12]), .C1(n29919), .O(n29920) );
  MAO222S U15533 ( .A1(n29931), .B1(rgb_value[11]), .C1(n29918), .O(n29919) );
  MAO222S U15534 ( .A1(n29933), .B1(rgb_value[10]), .C1(n29917), .O(n29918) );
  MAO222S U15535 ( .A1(rgb_value[8]), .B1(rgb_value[9]), .C1(n29936), .O(
        n29917) );
  MAO222 U15536 ( .A1(rgb_value[3]), .B1(n29949), .C1(n29938), .O(n29939) );
  MAO222S U15537 ( .A1(n29947), .B1(rgb_value[2]), .C1(n29937), .O(n29938) );
  MAO222S U15538 ( .A1(rgb_value[1]), .B1(rgb_value[0]), .C1(n29945), .O(
        n29937) );
  AO12S U15539 ( .B1(n24659), .B2(n24665), .A1(n24682), .O(n29312) );
  NR2 U15540 ( .I1(n24210), .I2(n24319), .O(n29227) );
  NR2 U15541 ( .I1(n24757), .I2(n24957), .O(n29392) );
  NR2 U15542 ( .I1(n24213), .I2(n24957), .O(n29280) );
  OA12S U15543 ( .B1(n24622), .B2(n24669), .A1(n24668), .O(n29364) );
  OA12S U15544 ( .B1(n24622), .B2(n24726), .A1(n24725), .O(n29351) );
  OA12S U15545 ( .B1(n24346), .B2(n24669), .A1(n24668), .O(n29273) );
  OA12S U15546 ( .B1(n24346), .B2(n24726), .A1(n24725), .O(n29267) );
  OA12S U15547 ( .B1(n24350), .B2(n24726), .A1(n24725), .O(n29264) );
  OA12S U15548 ( .B1(n24134), .B2(n24726), .A1(n24725), .O(n28629) );
  OA12 U15549 ( .B1(n24614), .B2(n24487), .A1(n24725), .O(n29070) );
  OA12 U15550 ( .B1(n24614), .B2(n23962), .A1(n24725), .O(n28626) );
  OA12 U15551 ( .B1(n24614), .B2(n24613), .A1(n24725), .O(n29355) );
  OA12S U15552 ( .B1(n24479), .B2(n24023), .A1(n24495), .O(n29054) );
  ND2 U15553 ( .I1(n24633), .I2(n24148), .O(n29207) );
  OA12 U15554 ( .B1(n24238), .B2(n24563), .A1(n24758), .O(n28672) );
  OA12 U15555 ( .B1(n24479), .B2(n24612), .A1(n24694), .O(n29233) );
  OA12S U15556 ( .B1(n24727), .B2(n24726), .A1(n24725), .O(n29405) );
  AO12S U15557 ( .B1(n24722), .B2(n24721), .A1(n24229), .O(n29402) );
  OA12 U15558 ( .B1(n24293), .B2(n24563), .A1(n24758), .O(n28729) );
  OA12 U15559 ( .B1(n24266), .B2(n24105), .A1(n24748), .O(n28722) );
  OA12S U15560 ( .B1(n24479), .B2(n24105), .A1(n24748), .O(n28612) );
  NR2 U15561 ( .I1(n24367), .I2(n24440), .O(n28821) );
  NR2 U15562 ( .I1(n24429), .I2(n24957), .O(n28804) );
  OA12S U15563 ( .B1(n24444), .B2(n24669), .A1(n24668), .O(n28857) );
  OA12S U15564 ( .B1(n24444), .B2(n24726), .A1(n24725), .O(n28845) );
  OA12S U15565 ( .B1(n24398), .B2(n24726), .A1(n24725), .O(n28848) );
  OA12S U15566 ( .B1(n24335), .B2(n24023), .A1(n24495), .O(n28778) );
  OA12S U15567 ( .B1(n24293), .B2(n24023), .A1(n24495), .O(n28736) );
  OA12 U15568 ( .B1(n24546), .B2(n24563), .A1(n24758), .O(n29115) );
  OA12S U15569 ( .B1(n24542), .B2(n24669), .A1(n24668), .O(n29084) );
  NR2 U15570 ( .I1(n24081), .I2(n24289), .O(n28740) );
  OA12S U15571 ( .B1(n24670), .B2(n24726), .A1(n24725), .O(n29309) );
  OA12S U15572 ( .B1(n24670), .B2(n24669), .A1(n24668), .O(n29321) );
  NR2 U15573 ( .I1(n24088), .I2(n24289), .O(n28747) );
  NR2 U15574 ( .I1(n24290), .I2(n24289), .O(n28969) );
  OA12S U15575 ( .B1(n24585), .B2(n24669), .A1(n24668), .O(n29163) );
  OA12S U15576 ( .B1(n24568), .B2(n24726), .A1(n24725), .O(n29148) );
  OA12S U15577 ( .B1(n24585), .B2(n24726), .A1(n24725), .O(n29151) );
  AO12S U15578 ( .B1(n24543), .B2(n24670), .A1(n24541), .O(n28761) );
  AO12 U15579 ( .B1(n24277), .B2(n24542), .A1(n24263), .O(n28712) );
  AO12 U15580 ( .B1(n24463), .B2(n24134), .A1(n24462), .O(n28602) );
  INV1 U15581 ( .I(n20769), .O(n29493) );
  AN2S U15582 ( .I1(n21389), .I2(n21388), .O(n13934) );
  ND2S U15583 ( .I1(n29521), .I2(n21619), .O(n21620) );
  ND2S U15584 ( .I1(n23107), .I2(n23100), .O(n23102) );
  ND2S U15585 ( .I1(n23098), .I2(n23097), .O(n23105) );
  ND2S U15586 ( .I1(n23096), .I2(n23095), .O(n23115) );
  ND2S U15587 ( .I1(n23034), .I2(n23033), .O(n23143) );
  ND2S U15588 ( .I1(n23025), .I2(n23024), .O(n23147) );
  ND2S U15589 ( .I1(n23011), .I2(n23010), .O(n23152) );
  ND2S U15590 ( .I1(n23008), .I2(n23007), .O(n23156) );
  ND2S U15591 ( .I1(n23006), .I2(n23005), .O(n23161) );
  OR2S U15592 ( .I1(n23002), .I2(n23003), .O(n23166) );
  OR2S U15593 ( .I1(n22831), .I2(n22832), .O(n22849) );
  ND2S U15594 ( .I1(n22830), .I2(n22829), .O(n22853) );
  OR2S U15595 ( .I1(n22829), .I2(n22830), .O(n22854) );
  ND2S U15596 ( .I1(n22806), .I2(n22805), .O(n22865) );
  ND2S U15597 ( .I1(n22762), .I2(n22761), .O(n22881) );
  ND2S U15598 ( .I1(n22753), .I2(n22752), .O(n22885) );
  ND2S U15599 ( .I1(n22739), .I2(n22738), .O(n22890) );
  ND2S U15600 ( .I1(n22736), .I2(n22735), .O(n22894) );
  HA1S U15601 ( .A(n22729), .B(n22728), .C(n22725), .S(n22903) );
  ND2S U15602 ( .I1(n23352), .I2(n23351), .O(n23368) );
  ND2S U15603 ( .I1(n23281), .I2(n23280), .O(n23401) );
  ND2S U15604 ( .I1(n23272), .I2(n23271), .O(n23405) );
  ND2S U15605 ( .I1(n23258), .I2(n23257), .O(n23410) );
  ND2S U15606 ( .I1(n23255), .I2(n23254), .O(n23414) );
  OR2S U15607 ( .I1(n23249), .I2(n23250), .O(n23424) );
  HA1 U15608 ( .A(n15988), .B(n15987), .C(n15989), .S(n23553) );
  ND2S U15609 ( .I1(n22589), .I2(n22582), .O(n22584) );
  ND2S U15610 ( .I1(n22580), .I2(n22579), .O(n22587) );
  ND2S U15611 ( .I1(n22503), .I2(n22502), .O(n22629) );
  ND2S U15612 ( .I1(n22489), .I2(n22488), .O(n22634) );
  ND2S U15613 ( .I1(n22486), .I2(n22485), .O(n22638) );
  ND2S U15614 ( .I1(n22484), .I2(n22483), .O(n22643) );
  OR2S U15615 ( .I1(n22480), .I2(n22481), .O(n22648) );
  ND2S U15616 ( .I1(n21979), .I2(n21972), .O(n21974) );
  ND2S U15617 ( .I1(n21970), .I2(n21969), .O(n21977) );
  ND2S U15618 ( .I1(n21905), .I2(n21904), .O(n22010) );
  ND2S U15619 ( .I1(n21903), .I2(n21902), .O(n22015) );
  ND2S U15620 ( .I1(n21894), .I2(n21893), .O(n22019) );
  ND2S U15621 ( .I1(n21880), .I2(n21879), .O(n22024) );
  ND2S U15622 ( .I1(n21877), .I2(n21876), .O(n22028) );
  ND2S U15623 ( .I1(n22231), .I2(n22224), .O(n22226) );
  ND2S U15624 ( .I1(n22222), .I2(n22221), .O(n22229) );
  ND2S U15625 ( .I1(n22155), .I2(n22154), .O(n22267) );
  ND2S U15626 ( .I1(n22146), .I2(n22145), .O(n22271) );
  ND2S U15627 ( .I1(n22132), .I2(n22131), .O(n22276) );
  ND2S U15628 ( .I1(n22129), .I2(n22128), .O(n22280) );
  ND2S U15629 ( .I1(n22127), .I2(n22126), .O(n22285) );
  OR2S U15630 ( .I1(n22123), .I2(n22124), .O(n22290) );
  ND2S U15631 ( .I1(n24031), .I2(n30004), .O(n13954) );
  ND2S U15632 ( .I1(n24701), .I2(n13950), .O(n13953) );
  ND2S U15633 ( .I1(addr[5]), .I2(addr[4]), .O(n23560) );
  ND2S U15634 ( .I1(n29552), .I2(n29549), .O(n29540) );
  ND2S U15635 ( .I1(n29552), .I2(n29547), .O(n29538) );
  ND2S U15636 ( .I1(col[0]), .I2(col[1]), .O(n24147) );
  ND3S U15637 ( .I1(n23651), .I2(n23649), .I3(n29964), .O(n23578) );
  AN2S U15638 ( .I1(action[1]), .I2(in_valid2), .O(n23654) );
  AN2S U15639 ( .I1(action[2]), .I2(in_valid2), .O(n23655) );
  AN2S U15640 ( .I1(action[0]), .I2(in_valid2), .O(n23663) );
  AN2S U15641 ( .I1(n29962), .I2(n23635), .O(n29961) );
  ND3S U15642 ( .I1(in_valid), .I2(n23690), .I3(n30005), .O(n30019) );
  ND2S U15643 ( .I1(set_cnt[1]), .I2(n29995), .O(n29997) );
  ND2S U15644 ( .I1(n30028), .I2(n23675), .O(n29999) );
  ND2S U15645 ( .I1(n13820), .I2(img[1912]), .O(n27945) );
  ND2S U15646 ( .I1(n13820), .I2(img[1914]), .O(n25772) );
  ND2S U15647 ( .I1(n13770), .I2(img[1272]), .O(n27925) );
  ND2S U15648 ( .I1(n13905), .I2(img[1392]), .O(n28294) );
  ND2S U15649 ( .I1(n13820), .I2(img[1394]), .O(n25441) );
  MUX2S U15650 ( .A(n28351), .B(img[544]), .S(n29481), .O(n12988) );
  MUX2S U15651 ( .A(n26826), .B(img[545]), .S(n29481), .O(n12987) );
  MUX2S U15652 ( .A(n29459), .B(img[547]), .S(n29481), .O(n12981) );
  MUX2S U15653 ( .A(n29337), .B(img[548]), .S(n29481), .O(n12982) );
  MUX2S U15654 ( .A(n29482), .B(img[549]), .S(n29481), .O(n12983) );
  MUX2S U15655 ( .A(n25214), .B(img[550]), .S(n29481), .O(n12984) );
  MUX2S U15656 ( .A(n24598), .B(img[551]), .S(n29481), .O(n12985) );
  MUX2S U15657 ( .A(n25781), .B(img[1698]), .S(n28922), .O(n11834) );
  MUX2S U15658 ( .A(n27620), .B(img[1955]), .S(n28993), .O(n11577) );
  MUX2S U15659 ( .A(n27146), .B(img[753]), .S(n29334), .O(n12779) );
  MUX2S U15660 ( .A(n29205), .B(img[740]), .S(n29204), .O(n12792) );
  MUX2S U15661 ( .A(n26105), .B(img[741]), .S(n29204), .O(n12791) );
  MUX2S U15662 ( .A(n24215), .B(img[743]), .S(n29204), .O(n12789) );
  MUX2S U15663 ( .A(n28459), .B(img[720]), .S(n29176), .O(n12812) );
  MUX2S U15664 ( .A(n28887), .B(img[708]), .S(n28886), .O(n12824) );
  MUX2S U15665 ( .A(n28002), .B(img[696]), .S(n28889), .O(n12836) );
  MUX2S U15666 ( .A(n27228), .B(img[697]), .S(n28889), .O(n12829) );
  MUX2S U15667 ( .A(n26008), .B(img[698]), .S(n28889), .O(n12830) );
  MUX2S U15668 ( .A(n27543), .B(img[699]), .S(n28889), .O(n12831) );
  MUX2S U15669 ( .A(n26428), .B(img[701]), .S(n28889), .O(n12833) );
  MUX2S U15670 ( .A(n24855), .B(img[702]), .S(n28889), .O(n12834) );
  MUX2S U15671 ( .A(n24427), .B(img[703]), .S(n28889), .O(n12835) );
  MUX2S U15672 ( .A(n28491), .B(img[688]), .S(n28666), .O(n12844) );
  MUX2S U15673 ( .A(n27192), .B(img[689]), .S(n28666), .O(n12843) );
  MUX2S U15674 ( .A(n25870), .B(img[690]), .S(n28666), .O(n12842) );
  MUX2S U15675 ( .A(n27739), .B(img[691]), .S(n28666), .O(n12841) );
  MUX2S U15676 ( .A(n28667), .B(img[692]), .S(n28666), .O(n12840) );
  MUX2S U15677 ( .A(n26479), .B(img[693]), .S(n28666), .O(n12839) );
  MUX2S U15678 ( .A(n25210), .B(img[694]), .S(n28666), .O(n12838) );
  MUX2S U15679 ( .A(n24004), .B(img[695]), .S(n28666), .O(n12837) );
  MUX2S U15680 ( .A(img[1804]), .B(n28687), .S(n28686), .O(n11728) );
  MUX2S U15681 ( .A(img[1548]), .B(n28744), .S(n28743), .O(n11984) );
  MUX2S U15682 ( .A(img[140]), .B(n29307), .S(n29306), .O(n13392) );
  MUX2S U15683 ( .A(img[372]), .B(n29316), .S(n29315), .O(n13160) );
  MUX2S U15684 ( .A(img[332]), .B(n28636), .S(n28635), .O(n13200) );
  MUX2S U15685 ( .A(img[316]), .B(n28855), .S(n28854), .O(n13216) );
  MUX2S U15686 ( .A(img[292]), .B(n29362), .S(n29361), .O(n13240) );
  MUX2S U15687 ( .A(img[908]), .B(n29301), .S(n29300), .O(n12624) );
  MUX2S U15688 ( .A(img[780]), .B(n29325), .S(n29324), .O(n12752) );
  MUX2S U15689 ( .A(img[652]), .B(n29332), .S(n29331), .O(n12880) );
  MUX2S U15690 ( .A(img[524]), .B(n29290), .S(n29289), .O(n13008) );
  MUX2S U15691 ( .A(img[1340]), .B(n28836), .S(n28835), .O(n12192) );
  MUX2S U15692 ( .A(img[1084]), .B(n28991), .S(n28990), .O(n12448) );
  MUX2S U15693 ( .A(img[1468]), .B(n28876), .S(n28875), .O(n12064) );
  MUX2S U15694 ( .A(img[956]), .B(n28843), .S(n28842), .O(n12576) );
  MUX2S U15695 ( .A(img[1460]), .B(n28653), .S(n28652), .O(n12072) );
  MUX2S U15696 ( .A(img[1204]), .B(n28599), .S(n28598), .O(n12328) );
  MUX2S U15697 ( .A(img[44]), .B(n29137), .S(n29136), .O(n13488) );
  MUX2S U15698 ( .A(img[1796]), .B(n28907), .S(n28906), .O(n11736) );
  MUX2S U15699 ( .A(img[1668]), .B(n28937), .S(n28936), .O(n11864) );
  MUX2S U15700 ( .A(img[1540]), .B(n28966), .S(n28965), .O(n11992) );
  MUX2S U15701 ( .A(img[1028]), .B(n28980), .S(n28979), .O(n12504) );
  MUX2S U15702 ( .A(img[772]), .B(n29424), .S(n29423), .O(n12760) );
  MUX2S U15703 ( .A(img[644]), .B(n29431), .S(n29430), .O(n12888) );
  MUX2S U15704 ( .A(img[260]), .B(n29410), .S(n29409), .O(n13272) );
  MUX2S U15705 ( .A(img[1020]), .B(n29400), .S(n29399), .O(n12512) );
  MUX2S U15706 ( .A(n29296), .B(img[12]), .S(n29295), .O(n13520) );
  MUX2S U15707 ( .A(n28642), .B(img[460]), .S(n28641), .O(n13072) );
  MUX2S U15708 ( .A(n29349), .B(img[932]), .S(n29348), .O(n12600) );
  MUX2S U15709 ( .A(n29375), .B(img[804]), .S(n29374), .O(n12728) );
  MUX2S U15710 ( .A(n29381), .B(img[676]), .S(n29380), .O(n12856) );
  MUX2S U15711 ( .A(n28772), .B(img[1964]), .S(n28771), .O(n11568) );
  MUX2S U15712 ( .A(n28702), .B(img[1708]), .S(n28701), .O(n11824) );
  MUX2S U15713 ( .A(n29390), .B(img[4]), .S(n29389), .O(n13528) );
  MUX2S U15714 ( .A(n29174), .B(img[684]), .S(n29173), .O(n12848) );
  MUX2S U15715 ( .A(n29231), .B(img[868]), .S(n29230), .O(n12664) );
  MUX2S U15716 ( .A(n28621), .B(img[948]), .S(n28620), .O(n12584) );
  MUX2S U15717 ( .A(n28660), .B(img[820]), .S(n28659), .O(n12712) );
  MUX2S U15718 ( .A(n28751), .B(img[1588]), .S(n28750), .O(n11944) );
  MUX2S U15719 ( .A(n29417), .B(img[388]), .S(n29416), .O(n13144) );
  MUX2S U15720 ( .A(img[407]), .B(n24502), .S(n29081), .O(n13125) );
  MUX2S U15721 ( .A(img[1807]), .B(n24039), .S(n28686), .O(n11725) );
  MUX2S U15722 ( .A(img[1551]), .B(n24085), .S(n28743), .O(n11981) );
  MUX2S U15723 ( .A(img[1295]), .B(n23940), .S(n28605), .O(n12237) );
  MUX2S U15724 ( .A(img[143]), .B(n24654), .S(n29306), .O(n13395) );
  MUX2S U15725 ( .A(img[663]), .B(n24533), .S(n29109), .O(n12869) );
  MUX2S U15726 ( .A(img[375]), .B(n24662), .S(n29315), .O(n13163) );
  MUX2S U15727 ( .A(img[343]), .B(n24561), .S(n29157), .O(n13195) );
  MUX2S U15728 ( .A(img[335]), .B(n23971), .S(n28635), .O(n13197) );
  MUX2S U15729 ( .A(img[295]), .B(n24593), .S(n29361), .O(n13243) );
  MUX2S U15730 ( .A(img[287]), .B(n24185), .S(n29179), .O(n13245) );
  MUX2S U15731 ( .A(img[911]), .B(n24648), .S(n29300), .O(n12627) );
  MUX2S U15732 ( .A(img[655]), .B(n24684), .S(n29331), .O(n12883) );
  MUX2S U15733 ( .A(img[527]), .B(n24642), .S(n29289), .O(n13005) );
  MUX2S U15734 ( .A(img[1599]), .B(n24281), .S(n28976), .O(n11933) );
  MUX2S U15735 ( .A(img[1087]), .B(n24441), .S(n28990), .O(n12445) );
  MUX2S U15736 ( .A(img[1463]), .B(n23990), .S(n28652), .O(n12069) );
  MUX2S U15737 ( .A(img[1207]), .B(n23934), .S(n28598), .O(n12325) );
  MUX2S U15738 ( .A(img[1799]), .B(n24230), .S(n28906), .O(n11739) );
  MUX2S U15739 ( .A(img[1671]), .B(n24260), .S(n28936), .O(n11861) );
  MUX2S U15740 ( .A(img[1543]), .B(n24286), .S(n28965), .O(n11995) );
  MUX2S U15741 ( .A(img[647]), .B(n24754), .S(n29430), .O(n12885) );
  MUX2S U15742 ( .A(img[263]), .B(n24730), .S(n29409), .O(n13275) );
  MUX2S U15743 ( .A(img[1023]), .B(n24719), .S(n29399), .O(n12515) );
  MUX2S U15744 ( .A(img[1183]), .B(n24160), .S(n29214), .O(n12355) );
  MUX2S U15745 ( .A(img[927]), .B(n24176), .S(n29221), .O(n12611) );
  MUX2S U15746 ( .A(img[543]), .B(n24141), .S(n29283), .O(n12989) );
  MUX2S U15747 ( .A(img[1055]), .B(n24320), .S(n29192), .O(n12477) );
  MUX2S U15748 ( .A(img[87]), .B(n24553), .S(n29139), .O(n13451) );
  MUX2S U15749 ( .A(img[79]), .B(n23912), .S(n28587), .O(n13453) );
  MUX2S U15750 ( .A(img[31]), .B(n24145), .S(n29276), .O(n13501) );
  MUX2S U15751 ( .A(img[1679]), .B(n24063), .S(n28715), .O(n11859) );
  MUX2S U15752 ( .A(img[1039]), .B(n24100), .S(n28757), .O(n12493) );
  MUX2S U15753 ( .A(n24767), .B(img[15]), .S(n29295), .O(n13517) );
  MUX2S U15754 ( .A(n23980), .B(img[463]), .S(n28641), .O(n13075) );
  MUX2S U15755 ( .A(n24607), .B(img[935]), .S(n29348), .O(n12597) );
  MUX2S U15756 ( .A(n24634), .B(img[679]), .S(n29380), .O(n12853) );
  MUX2S U15757 ( .A(n24114), .B(img[1967]), .S(n28771), .O(n11571) );
  MUX2S U15758 ( .A(n24053), .B(img[1711]), .S(n28701), .O(n11827) );
  MUX2S U15759 ( .A(n24709), .B(img[7]), .S(n29389), .O(n13525) );
  MUX2S U15760 ( .A(n24591), .B(img[943]), .S(n29142), .O(n12589) );
  MUX2S U15761 ( .A(n24583), .B(img[687]), .S(n29173), .O(n12851) );
  MUX2S U15762 ( .A(n24131), .B(img[1975]), .S(n28792), .O(n11557) );
  MUX2S U15763 ( .A(n23952), .B(img[951]), .S(n28620), .O(n12581) );
  MUX2S U15764 ( .A(img[529]), .B(n27232), .S(n29021), .O(n12997) );
  MUX2S U15765 ( .A(img[534]), .B(n25358), .S(n29021), .O(n13002) );
  MUX2S U15766 ( .A(img[401]), .B(n27252), .S(n29081), .O(n13131) );
  MUX2S U15767 ( .A(img[406]), .B(n25379), .S(n29081), .O(n13126) );
  MUX2S U15768 ( .A(n24690), .B(img[519]), .S(n29383), .O(n13019) );
  MUX2S U15769 ( .A(img[1806]), .B(n25031), .S(n28686), .O(n11726) );
  MUX2S U15770 ( .A(img[1550]), .B(n25072), .S(n28743), .O(n11982) );
  MUX2S U15771 ( .A(img[1294]), .B(n24976), .S(n28605), .O(n12238) );
  MUX2S U15772 ( .A(img[137]), .B(n27122), .S(n29306), .O(n13389) );
  MUX2S U15773 ( .A(img[142]), .B(n24985), .S(n29306), .O(n13394) );
  MUX2S U15774 ( .A(img[657]), .B(n27261), .S(n29109), .O(n12875) );
  MUX2S U15775 ( .A(img[662]), .B(n25388), .S(n29109), .O(n12870) );
  MUX2S U15776 ( .A(img[369]), .B(n27128), .S(n29315), .O(n13157) );
  MUX2S U15777 ( .A(img[374]), .B(n24991), .S(n29315), .O(n13162) );
  MUX2S U15778 ( .A(img[329]), .B(n27182), .S(n28635), .O(n13203) );
  MUX2S U15779 ( .A(img[313]), .B(n27214), .S(n28854), .O(n13219) );
  MUX2S U15780 ( .A(img[318]), .B(n24831), .S(n28854), .O(n13214) );
  MUX2S U15781 ( .A(img[302]), .B(n25343), .S(n29154), .O(n13230) );
  MUX2S U15782 ( .A(img[289]), .B(n26863), .S(n29361), .O(n13237) );
  MUX2S U15783 ( .A(img[294]), .B(n25230), .S(n29361), .O(n13242) );
  MUX2S U15784 ( .A(img[281]), .B(n26916), .S(n29179), .O(n13251) );
  MUX2S U15785 ( .A(img[1161]), .B(n27093), .S(n28590), .O(n12365) );
  MUX2S U15786 ( .A(img[1166]), .B(n24966), .S(n28590), .O(n12370) );
  MUX2S U15787 ( .A(img[654]), .B(n25012), .S(n29331), .O(n12882) );
  MUX2S U15788 ( .A(img[521]), .B(n27103), .S(n29289), .O(n13011) );
  MUX2S U15789 ( .A(img[526]), .B(n24951), .S(n29289), .O(n13006) );
  MUX2S U15790 ( .A(n24046), .B(img[1847]), .S(n28693), .O(n11691) );
  MUX2S U15791 ( .A(n24666), .B(img[399]), .S(n29318), .O(n13139) );
  MUX2S U15792 ( .A(n24058), .B(img[1687]), .S(n28708), .O(n11845) );
  MUX2S U15793 ( .A(img[1726]), .B(n24895), .S(n28948), .O(n11810) );
  MUX2S U15794 ( .A(img[1337]), .B(n26690), .S(n28835), .O(n12195) );
  MUX2S U15795 ( .A(img[1342]), .B(n24818), .S(n28835), .O(n12190) );
  MUX2S U15796 ( .A(img[1081]), .B(n26795), .S(n28990), .O(n12451) );
  MUX2S U15797 ( .A(img[1465]), .B(n26717), .S(n28875), .O(n12061) );
  MUX2S U15798 ( .A(img[273]), .B(n27248), .S(n29074), .O(n13253) );
  MUX2S U15799 ( .A(img[278]), .B(n25374), .S(n29074), .O(n13258) );
  MUX2S U15800 ( .A(img[1457]), .B(n27134), .S(n28652), .O(n12075) );
  MUX2S U15801 ( .A(img[1462]), .B(n24997), .S(n28652), .O(n12070) );
  MUX2S U15802 ( .A(img[1201]), .B(n27088), .S(n28598), .O(n12331) );
  MUX2S U15803 ( .A(img[1206]), .B(n24961), .S(n28598), .O(n12326) );
  MUX2S U15804 ( .A(img[1793]), .B(n26753), .S(n28906), .O(n11733) );
  MUX2S U15805 ( .A(img[1665]), .B(n26773), .S(n28936), .O(n11867) );
  MUX2S U15806 ( .A(img[1670]), .B(n24889), .S(n28936), .O(n11862) );
  MUX2S U15807 ( .A(img[1537]), .B(n26793), .S(n28965), .O(n11989) );
  MUX2S U15808 ( .A(img[1542]), .B(n24910), .S(n28965), .O(n11994) );
  MUX2S U15809 ( .A(img[1414]), .B(n24839), .S(n28864), .O(n12118) );
  MUX2S U15810 ( .A(img[1281]), .B(n26698), .S(n28824), .O(n12245) );
  MUX2S U15811 ( .A(img[1158]), .B(n24802), .S(n28810), .O(n12374) );
  MUX2S U15812 ( .A(img[1030]), .B(n24920), .S(n28979), .O(n12506) );
  MUX2S U15813 ( .A(img[641]), .B(n26733), .S(n29430), .O(n12891) );
  MUX2S U15814 ( .A(img[646]), .B(n25278), .S(n29430), .O(n12886) );
  MUX2S U15815 ( .A(img[257]), .B(n26710), .S(n29409), .O(n13269) );
  MUX2S U15816 ( .A(img[262]), .B(n25252), .S(n29409), .O(n13274) );
  MUX2S U15817 ( .A(img[1430]), .B(n25292), .S(n29094), .O(n12102) );
  MUX2S U15818 ( .A(img[1174]), .B(n25321), .S(n29040), .O(n12358) );
  MUX2S U15819 ( .A(img[1017]), .B(n26700), .S(n29399), .O(n12509) );
  MUX2S U15820 ( .A(img[1022]), .B(n25267), .S(n29399), .O(n12514) );
  MUX2S U15821 ( .A(img[1009]), .B(n27161), .S(n29303), .O(n12523) );
  MUX2S U15822 ( .A(img[1014]), .B(n24983), .S(n29303), .O(n12518) );
  MUX2S U15823 ( .A(img[1001]), .B(n27238), .S(n29064), .O(n12525) );
  MUX2S U15824 ( .A(img[1006]), .B(n25368), .S(n29064), .O(n12530) );
  MUX2S U15825 ( .A(img[961]), .B(n27204), .S(n28838), .O(n12571) );
  MUX2S U15826 ( .A(img[966]), .B(n24825), .S(n28838), .O(n12566) );
  MUX2S U15827 ( .A(img[1193]), .B(n26944), .S(n29033), .O(n12333) );
  MUX2S U15828 ( .A(img[1177]), .B(n26832), .S(n29214), .O(n12349) );
  MUX2S U15829 ( .A(img[921]), .B(n26908), .S(n29221), .O(n12605) );
  MUX2S U15830 ( .A(img[665]), .B(n26929), .S(n29201), .O(n12861) );
  MUX2S U15831 ( .A(img[537]), .B(n26900), .S(n29283), .O(n12995) );
  MUX2S U15832 ( .A(img[105]), .B(n27234), .S(n29030), .O(n13427) );
  MUX2S U15833 ( .A(img[110]), .B(n25364), .S(n29030), .O(n13422) );
  MUX2S U15834 ( .A(img[1822]), .B(n24864), .S(n28899), .O(n11710) );
  MUX2S U15835 ( .A(img[1561]), .B(n26780), .S(n28958), .O(n11971) );
  MUX2S U15836 ( .A(img[1566]), .B(n24905), .S(n28958), .O(n11966) );
  MUX2S U15837 ( .A(img[1049]), .B(n26888), .S(n29192), .O(n12483) );
  MUX2S U15838 ( .A(img[409]), .B(n26920), .S(n29270), .O(n13117) );
  MUX2S U15839 ( .A(img[81]), .B(n26937), .S(n29139), .O(n13445) );
  MUX2S U15840 ( .A(img[86]), .B(n25317), .S(n29139), .O(n13450) );
  MUX2S U15841 ( .A(img[73]), .B(n27169), .S(n28587), .O(n13459) );
  MUX2S U15842 ( .A(img[57]), .B(n27202), .S(n28807), .O(n13475) );
  MUX2S U15843 ( .A(img[62]), .B(n24798), .S(n28807), .O(n13470) );
  MUX2S U15844 ( .A(img[33]), .B(n26830), .S(n29342), .O(n13493) );
  MUX2S U15845 ( .A(img[25]), .B(n26904), .S(n29276), .O(n13507) );
  MUX2S U15846 ( .A(img[441]), .B(n27218), .S(n28860), .O(n13086) );
  MUX2S U15847 ( .A(img[446]), .B(n24835), .S(n28860), .O(n13091) );
  MUX2S U15848 ( .A(img[150]), .B(n25370), .S(n29067), .O(n13382) );
  MUX2S U15849 ( .A(img[1689]), .B(n26760), .S(n28929), .O(n11837) );
  MUX2S U15850 ( .A(img[1694]), .B(n24884), .S(n28929), .O(n11842) );
  MUX2S U15851 ( .A(img[1678]), .B(n25051), .S(n28715), .O(n11858) );
  MUX2S U15852 ( .A(img[1033]), .B(n27153), .S(n28757), .O(n12499) );
  MUX2S U15853 ( .A(img[1038]), .B(n25082), .S(n28757), .O(n12494) );
  MUX2S U15854 ( .A(n24955), .B(img[14]), .S(n29295), .O(n13518) );
  MUX2S U15855 ( .A(n27184), .B(img[433]), .S(n28638), .O(n13099) );
  MUX2S U15856 ( .A(n25201), .B(img[438]), .S(n28638), .O(n13094) );
  MUX2S U15857 ( .A(n26854), .B(img[929]), .S(n29348), .O(n12603) );
  MUX2S U15858 ( .A(n26886), .B(img[673]), .S(n29380), .O(n12859) );
  MUX2S U15859 ( .A(n25243), .B(img[678]), .S(n29380), .O(n12854) );
  MUX2S U15860 ( .A(n25036), .B(img[1710]), .S(n28701), .O(n11826) );
  MUX2S U15861 ( .A(n26678), .B(img[1]), .S(n29389), .O(n13531) );
  MUX2S U15862 ( .A(n25261), .B(img[6]), .S(n29389), .O(n13526) );
  MUX2S U15863 ( .A(n25334), .B(img[942]), .S(n29142), .O(n12590) );
  MUX2S U15864 ( .A(n25356), .B(img[686]), .S(n29173), .O(n12850) );
  MUX2S U15865 ( .A(n26727), .B(img[889]), .S(n29427), .O(n12643) );
  MUX2S U15866 ( .A(n27190), .B(img[841]), .S(n28663), .O(n12691) );
  MUX2S U15867 ( .A(n27172), .B(img[945]), .S(n28620), .O(n12587) );
  MUX2S U15868 ( .A(n25067), .B(img[1590]), .S(n28750), .O(n11946) );
  MUX2S U15869 ( .A(n26674), .B(img[513]), .S(n29383), .O(n13013) );
  MUX2S U15870 ( .A(n25256), .B(img[518]), .S(n29383), .O(n13018) );
  MUX2S U15871 ( .A(n28212), .B(img[1704]), .S(n28701), .O(n11828) );
  MUX2S U15872 ( .A(n27030), .B(img[1705]), .S(n28701), .O(n11821) );
  MUX2S U15873 ( .A(n25507), .B(img[1706]), .S(n28701), .O(n11822) );
  MUX2S U15874 ( .A(n26735), .B(img[1825]), .S(n28892), .O(n11701) );
  MUX2S U15875 ( .A(n27025), .B(img[1681]), .S(n28708), .O(n11851) );
  MUX2S U15876 ( .A(n25041), .B(img[1686]), .S(n28708), .O(n11846) );
  MUX2S U15877 ( .A(n28264), .B(img[1960]), .S(n28771), .O(n11572) );
  MUX2S U15878 ( .A(n27438), .B(img[1963]), .S(n28771), .O(n11567) );
  MUX2S U15879 ( .A(n26345), .B(img[1965]), .S(n28771), .O(n11569) );
  MUX2S U15880 ( .A(n28253), .B(img[1968]), .S(n28792), .O(n11564) );
  MUX2S U15881 ( .A(n27793), .B(img[931]), .S(n29348), .O(n12601) );
  MUX2S U15882 ( .A(n26615), .B(img[933]), .S(n29348), .O(n12599) );
  MUX2S U15883 ( .A(n25222), .B(img[934]), .S(n29348), .O(n12598) );
  MUX2S U15884 ( .A(n26991), .B(img[681]), .S(n29173), .O(n12845) );
  MUX2S U15885 ( .A(n25638), .B(img[682]), .S(n29173), .O(n12846) );
  MUX2S U15886 ( .A(n27480), .B(img[683]), .S(n29173), .O(n12847) );
  MUX2S U15887 ( .A(n26460), .B(img[685]), .S(n29173), .O(n12849) );
  MUX2S U15888 ( .A(img[528]), .B(n28116), .S(n29021), .O(n13004) );
  MUX2S U15889 ( .A(img[530]), .B(n25662), .S(n29021), .O(n12998) );
  MUX2S U15890 ( .A(img[400]), .B(n28157), .S(n29081), .O(n13132) );
  MUX2S U15891 ( .A(img[402]), .B(n25678), .S(n29081), .O(n13130) );
  MUX2S U15892 ( .A(img[1800]), .B(n28187), .S(n28686), .O(n11732) );
  MUX2S U15893 ( .A(img[1802]), .B(n25505), .S(n28686), .O(n11730) );
  MUX2S U15894 ( .A(img[1546]), .B(n25545), .S(n28743), .O(n11986) );
  MUX2S U15895 ( .A(img[1290]), .B(n25449), .S(n28605), .O(n12242) );
  MUX2S U15896 ( .A(img[656]), .B(n28177), .S(n29109), .O(n12876) );
  MUX2S U15897 ( .A(img[658]), .B(n25654), .S(n29109), .O(n12874) );
  MUX2S U15898 ( .A(img[370]), .B(n25459), .S(n29315), .O(n13158) );
  MUX2S U15899 ( .A(img[328]), .B(n28480), .S(n28635), .O(n13204) );
  MUX2S U15900 ( .A(img[330]), .B(n25868), .S(n28635), .O(n13202) );
  MUX2S U15901 ( .A(img[312]), .B(n27986), .S(n28854), .O(n13220) );
  MUX2S U15902 ( .A(img[314]), .B(n25994), .S(n28854), .O(n13218) );
  MUX2S U15903 ( .A(img[296]), .B(n28444), .S(n29154), .O(n13236) );
  MUX2S U15904 ( .A(img[298]), .B(n25615), .S(n29154), .O(n13234) );
  MUX2S U15905 ( .A(img[288]), .B(n28388), .S(n29361), .O(n13244) );
  MUX2S U15906 ( .A(img[290]), .B(n25902), .S(n29361), .O(n13238) );
  MUX2S U15907 ( .A(img[280]), .B(n28511), .S(n29179), .O(n13252) );
  MUX2S U15908 ( .A(img[282]), .B(n25966), .S(n29179), .O(n13250) );
  MUX2S U15909 ( .A(img[1162]), .B(n25438), .S(n28590), .O(n12366) );
  MUX2S U15910 ( .A(img[648]), .B(n28337), .S(n29331), .O(n12884) );
  MUX2S U15911 ( .A(img[650]), .B(n25485), .S(n29331), .O(n12878) );
  MUX2S U15912 ( .A(img[522]), .B(n25424), .S(n29289), .O(n13010) );
  MUX2S U15913 ( .A(img[1592]), .B(n28042), .S(n28976), .O(n11940) );
  MUX2S U15914 ( .A(img[1336]), .B(n27973), .S(n28835), .O(n12196) );
  MUX2S U15915 ( .A(img[1080]), .B(n28053), .S(n28990), .O(n12452) );
  MUX2S U15916 ( .A(img[1464]), .B(n27959), .S(n28875), .O(n12068) );
  MUX2S U15917 ( .A(img[272]), .B(n28153), .S(n29074), .O(n13260) );
  MUX2S U15918 ( .A(img[274]), .B(n25658), .S(n29074), .O(n13254) );
  MUX2S U15919 ( .A(img[1202]), .B(n25430), .S(n28598), .O(n12330) );
  MUX2S U15920 ( .A(img[1792]), .B(n27939), .S(n28906), .O(n11740) );
  MUX2S U15921 ( .A(img[1664]), .B(n28016), .S(n28936), .O(n11868) );
  MUX2S U15922 ( .A(img[1536]), .B(n28036), .S(n28965), .O(n11996) );
  MUX2S U15923 ( .A(img[1152]), .B(n27918), .S(n28810), .O(n12380) );
  MUX2S U15924 ( .A(img[1154]), .B(n25690), .S(n28810), .O(n12378) );
  MUX2S U15925 ( .A(img[640]), .B(n28114), .S(n29430), .O(n12892) );
  MUX2S U15926 ( .A(img[256]), .B(n28099), .S(n29409), .O(n13276) );
  MUX2S U15927 ( .A(img[1426]), .B(n25623), .S(n29094), .O(n12106) );
  MUX2S U15928 ( .A(img[1168]), .B(n28129), .S(n29040), .O(n12364) );
  MUX2S U15929 ( .A(img[1016]), .B(n28089), .S(n29399), .O(n12516) );
  MUX2S U15930 ( .A(img[1010]), .B(n25451), .S(n29303), .O(n12522) );
  MUX2S U15931 ( .A(img[1000]), .B(n28147), .S(n29064), .O(n12532) );
  MUX2S U15932 ( .A(img[1002]), .B(n25668), .S(n29064), .O(n12526) );
  MUX2S U15933 ( .A(img[984]), .B(n28381), .S(n29345), .O(n12548) );
  MUX2S U15934 ( .A(img[986]), .B(n25946), .S(n29345), .O(n12542) );
  MUX2S U15935 ( .A(img[960]), .B(n27980), .S(n28838), .O(n12572) );
  MUX2S U15936 ( .A(img[962]), .B(n25988), .S(n28838), .O(n12570) );
  MUX2S U15937 ( .A(img[1194]), .B(n25590), .S(n29033), .O(n12334) );
  MUX2S U15938 ( .A(img[1178]), .B(n25878), .S(n29214), .O(n12350) );
  MUX2S U15939 ( .A(img[920]), .B(n28503), .S(n29221), .O(n12612) );
  MUX2S U15940 ( .A(img[922]), .B(n25958), .S(n29221), .O(n12606) );
  MUX2S U15941 ( .A(img[664]), .B(n28524), .S(n29201), .O(n12868) );
  MUX2S U15942 ( .A(img[666]), .B(n25978), .S(n29201), .O(n12862) );
  MUX2S U15943 ( .A(img[536]), .B(n28495), .S(n29283), .O(n12996) );
  MUX2S U15944 ( .A(img[538]), .B(n25950), .S(n29283), .O(n12994) );
  MUX2S U15945 ( .A(img[104]), .B(n28122), .S(n29030), .O(n13428) );
  MUX2S U15946 ( .A(img[106]), .B(n25664), .S(n29030), .O(n13426) );
  MUX2S U15947 ( .A(img[114]), .B(n25426), .S(n29536), .O(n13414) );
  MUX2S U15948 ( .A(img[1816]), .B(n27934), .S(n28899), .O(n11716) );
  MUX2S U15949 ( .A(img[1048]), .B(n28417), .S(n29192), .O(n12484) );
  MUX2S U15950 ( .A(img[1050]), .B(n25930), .S(n29192), .O(n12482) );
  MUX2S U15951 ( .A(img[408]), .B(n28515), .S(n29270), .O(n13124) );
  MUX2S U15952 ( .A(img[410]), .B(n25970), .S(n29270), .O(n13118) );
  MUX2S U15953 ( .A(img[80]), .B(n28437), .S(n29139), .O(n13452) );
  MUX2S U15954 ( .A(img[82]), .B(n25583), .S(n29139), .O(n13446) );
  MUX2S U15955 ( .A(img[72]), .B(n28467), .S(n28587), .O(n13460) );
  MUX2S U15956 ( .A(img[74]), .B(n25846), .S(n28587), .O(n13458) );
  MUX2S U15957 ( .A(img[56]), .B(n27964), .S(n28807), .O(n13476) );
  MUX2S U15958 ( .A(img[58]), .B(n25982), .S(n28807), .O(n13474) );
  MUX2S U15959 ( .A(img[34]), .B(n25874), .S(n29342), .O(n13494) );
  MUX2S U15960 ( .A(img[24]), .B(n28499), .S(n29276), .O(n13508) );
  MUX2S U15961 ( .A(img[26]), .B(n25954), .S(n29276), .O(n13506) );
  MUX2S U15962 ( .A(img[440]), .B(n27992), .S(n28860), .O(n13092) );
  MUX2S U15963 ( .A(img[442]), .B(n25998), .S(n28860), .O(n13087) );
  MUX2S U15964 ( .A(img[424]), .B(n28448), .S(n29160), .O(n13108) );
  MUX2S U15965 ( .A(img[418]), .B(n25907), .S(n29367), .O(n13114) );
  MUX2S U15966 ( .A(img[1688]), .B(n28011), .S(n28929), .O(n11844) );
  MUX2S U15967 ( .A(img[1674]), .B(n25525), .S(n28715), .O(n11854) );
  MUX2S U15968 ( .A(img[1032]), .B(n28349), .S(n28757), .O(n12500) );
  MUX2S U15969 ( .A(img[1034]), .B(n25555), .S(n28757), .O(n12498) );
  MUX2S U15970 ( .A(n28482), .B(img[432]), .S(n28638), .O(n13100) );
  MUX2S U15971 ( .A(n25856), .B(img[434]), .S(n28638), .O(n13098) );
  MUX2S U15972 ( .A(n28411), .B(img[672]), .S(n29380), .O(n12860) );
  MUX2S U15973 ( .A(n25926), .B(img[674]), .S(n29380), .O(n12858) );
  MUX2S U15974 ( .A(n28422), .B(img[1056]), .S(n29185), .O(n12476) );
  MUX2S U15975 ( .A(n28087), .B(img[0]), .S(n29389), .O(n13532) );
  MUX2S U15976 ( .A(n25628), .B(img[1450]), .S(n29087), .O(n12078) );
  MUX2S U15977 ( .A(n28439), .B(img[936]), .S(n29142), .O(n12596) );
  MUX2S U15978 ( .A(n25607), .B(img[938]), .S(n29142), .O(n12592) );
  MUX2S U15979 ( .A(n25972), .B(img[866]), .S(n29230), .O(n12662) );
  MUX2S U15980 ( .A(n25602), .B(img[1322]), .S(n29047), .O(n12210) );
  MUX2S U15981 ( .A(n28470), .B(img[944]), .S(n28620), .O(n12588) );
  MUX2S U15982 ( .A(n25848), .B(img[946]), .S(n28620), .O(n12586) );
  MUX2S U15983 ( .A(n25537), .B(img[1586]), .S(n28750), .O(n11942) );
  MUX2S U15984 ( .A(n28082), .B(img[512]), .S(n29383), .O(n13020) );
  MUX2S U15985 ( .A(n27929), .B(img[1824]), .S(n28892), .O(n11708) );
  MUX2S U15986 ( .A(img[532]), .B(n29022), .S(n29021), .O(n13000) );
  MUX2S U15987 ( .A(img[404]), .B(n29082), .S(n29081), .O(n13128) );
  MUX2S U15988 ( .A(n25476), .B(img[1418]), .S(n28645), .O(n12110) );
  MUX2S U15989 ( .A(n28197), .B(img[1808]), .S(n28679), .O(n11724) );
  MUX2S U15990 ( .A(n25512), .B(img[1682]), .S(n28708), .O(n11850) );
  MUX2S U15991 ( .A(img[916]), .B(n29062), .S(n29061), .O(n12616) );
  MUX2S U15992 ( .A(img[788]), .B(n29103), .S(n29102), .O(n12744) );
  MUX2S U15993 ( .A(img[660]), .B(n29110), .S(n29109), .O(n12872) );
  MUX2S U15994 ( .A(img[20]), .B(n29028), .S(n29027), .O(n13512) );
  MUX2S U15995 ( .A(img[276]), .B(n29075), .S(n29074), .O(n13256) );
  MUX2S U15996 ( .A(img[1172]), .B(n29041), .S(n29040), .O(n12360) );
  MUX2S U15997 ( .A(n29088), .B(img[1452]), .S(n29087), .O(n12080) );
  MUX2S U15998 ( .A(n29048), .B(img[1324]), .S(n29047), .O(n12208) );
  MUX2S U15999 ( .A(img[319]), .B(n24394), .S(n28854), .O(n13213) );
  MUX2S U16000 ( .A(n29143), .B(img[940]), .S(n29142), .O(n12594) );
  MUX2S U16001 ( .A(n26440), .B(img[941]), .S(n29142), .O(n12595) );
  MUX2S U16002 ( .A(img[1471]), .B(n24410), .S(n28875), .O(n12067) );
  MUX2S U16003 ( .A(img[1415]), .B(n24403), .S(n28864), .O(n12117) );
  MUX2S U16004 ( .A(img[1287]), .B(n24373), .S(n28824), .O(n12251) );
  MUX2S U16005 ( .A(img[967]), .B(n24388), .S(n28838), .O(n12565) );
  MUX2S U16006 ( .A(img[63]), .B(n24358), .S(n28807), .O(n13469) );
  MUX2S U16007 ( .A(img[447]), .B(n24399), .S(n28860), .O(n13085) );
  MUX2S U16008 ( .A(img[531]), .B(n27293), .S(n29021), .O(n12999) );
  MUX2S U16009 ( .A(img[403]), .B(n27333), .S(n29081), .O(n13129) );
  MUX2S U16010 ( .A(img[1547]), .B(n27403), .S(n28743), .O(n11985) );
  MUX2S U16011 ( .A(img[659]), .B(n27352), .S(n29109), .O(n12873) );
  MUX2S U16012 ( .A(img[355]), .B(n27874), .S(n29182), .O(n13175) );
  MUX2S U16013 ( .A(img[331]), .B(n27732), .S(n28635), .O(n13201) );
  MUX2S U16014 ( .A(img[315]), .B(n27519), .S(n28854), .O(n13217) );
  MUX2S U16015 ( .A(img[299]), .B(n27468), .S(n29154), .O(n13233) );
  MUX2S U16016 ( .A(img[291]), .B(n27815), .S(n29361), .O(n13239) );
  MUX2S U16017 ( .A(img[1339]), .B(n27505), .S(n28835), .O(n12193) );
  MUX2S U16018 ( .A(img[19]), .B(n27297), .S(n29027), .O(n13511) );
  MUX2S U16019 ( .A(img[955]), .B(n27510), .S(n28842), .O(n12575) );
  MUX2S U16020 ( .A(img[275]), .B(n27329), .S(n29074), .O(n13255) );
  MUX2S U16021 ( .A(img[43]), .B(n27456), .S(n29136), .O(n13489) );
  MUX2S U16022 ( .A(img[1801]), .B(n27000), .S(n28686), .O(n11731) );
  MUX2S U16023 ( .A(img[297]), .B(n26967), .S(n29154), .O(n13235) );
  MUX2S U16024 ( .A(img[286]), .B(n25145), .S(n29179), .O(n13246) );
  MUX2S U16025 ( .A(img[1795]), .B(n27557), .S(n28906), .O(n11735) );
  MUX2S U16026 ( .A(img[1411]), .B(n27527), .S(n28864), .O(n12121) );
  MUX2S U16027 ( .A(img[899]), .B(n27835), .S(n29395), .O(n12633) );
  MUX2S U16028 ( .A(img[643]), .B(n27852), .S(n29430), .O(n12889) );
  MUX2S U16029 ( .A(img[259]), .B(n27843), .S(n29409), .O(n13271) );
  MUX2S U16030 ( .A(img[1427]), .B(n27344), .S(n29094), .O(n12105) );
  MUX2S U16031 ( .A(img[1171]), .B(n27307), .S(n29040), .O(n12361) );
  MUX2S U16032 ( .A(img[1003]), .B(n27319), .S(n29064), .O(n12527) );
  MUX2S U16033 ( .A(img[979]), .B(n27458), .S(n29145), .O(n12553) );
  MUX2S U16034 ( .A(img[923]), .B(n27864), .S(n29221), .O(n12607) );
  MUX2S U16035 ( .A(img[667]), .B(n27884), .S(n29201), .O(n12863) );
  MUX2S U16036 ( .A(img[539]), .B(n27856), .S(n29283), .O(n12993) );
  MUX2S U16037 ( .A(img[1051]), .B(n27756), .S(n29192), .O(n12481) );
  MUX2S U16038 ( .A(img[411]), .B(n27876), .S(n29270), .O(n13119) );
  MUX2S U16039 ( .A(img[35]), .B(n27768), .S(n29342), .O(n13495) );
  MUX2S U16040 ( .A(img[27]), .B(n27860), .S(n29276), .O(n13505) );
  MUX2S U16041 ( .A(img[427]), .B(n27472), .S(n29160), .O(n13103) );
  MUX2S U16042 ( .A(img[1675]), .B(n27383), .S(n28715), .O(n11855) );
  MUX2S U16043 ( .A(img[1035]), .B(n27715), .S(n28757), .O(n12497) );
  MUX2S U16044 ( .A(img[1425]), .B(n26976), .S(n29094), .O(n12107) );
  MUX2S U16045 ( .A(n27743), .B(img[435]), .S(n28638), .O(n13097) );
  MUX2S U16046 ( .A(img[977]), .B(n26961), .S(n29145), .O(n12555) );
  MUX2S U16047 ( .A(n27806), .B(img[1443]), .S(n29248), .O(n12089) );
  MUX2S U16048 ( .A(n27811), .B(img[675]), .S(n29380), .O(n12857) );
  MUX2S U16049 ( .A(img[926]), .B(n25137), .S(n29221), .O(n12610) );
  MUX2S U16050 ( .A(img[670]), .B(n25169), .S(n29201), .O(n12866) );
  MUX2S U16051 ( .A(img[542]), .B(n25109), .S(n29283), .O(n12990) );
  MUX2S U16052 ( .A(img[414]), .B(n25149), .S(n29270), .O(n13122) );
  MUX2S U16053 ( .A(img[30]), .B(n25113), .S(n29276), .O(n13502) );
  MUX2S U16054 ( .A(img[425]), .B(n26972), .S(n29160), .O(n13101) );
  MUX2S U16055 ( .A(img[1673]), .B(n27020), .S(n28715), .O(n11853) );
  MUX2S U16056 ( .A(n27831), .B(img[3]), .S(n29389), .O(n13529) );
  MUX2S U16057 ( .A(n27346), .B(img[875]), .S(n29106), .O(n12657) );
  MUX2S U16058 ( .A(n27882), .B(img[867]), .S(n29230), .O(n12663) );
  MUX2S U16059 ( .A(n27821), .B(img[859]), .S(n29371), .O(n12673) );
  MUX2S U16060 ( .A(n27474), .B(img[851]), .S(n29170), .O(n12679) );
  MUX2S U16061 ( .A(n27721), .B(img[947]), .S(n28620), .O(n12585) );
  MUX2S U16062 ( .A(n27734), .B(img[819]), .S(n28659), .O(n12711) );
  MUX2S U16063 ( .A(n27827), .B(img[515]), .S(n29383), .O(n13015) );
  MUX2S U16064 ( .A(n27823), .B(img[387]), .S(n29416), .O(n13145) );
  MUX2S U16065 ( .A(n27375), .B(img[1811]), .S(n28679), .O(n11719) );
  MUX2S U16066 ( .A(n27396), .B(img[1683]), .S(n28708), .O(n11849) );
  MUX2S U16067 ( .A(n27426), .B(img[1043]), .S(n29122), .O(n12486) );
  MUX2S U16068 ( .A(n26954), .B(img[1321]), .S(n29047), .O(n12211) );
  MUX2S U16069 ( .A(n28317), .B(img[392]), .S(n29318), .O(n13140) );
  MUX2S U16070 ( .A(n27684), .B(img[395]), .S(n29318), .O(n13135) );
  MUX2S U16071 ( .A(img[1805]), .B(n26269), .S(n28686), .O(n11727) );
  MUX2S U16072 ( .A(img[1544]), .B(n28228), .S(n28743), .O(n11988) );
  MUX2S U16073 ( .A(img[1545]), .B(n27040), .S(n28743), .O(n11987) );
  MUX2S U16074 ( .A(img[1549]), .B(n26309), .S(n28743), .O(n11983) );
  MUX2S U16075 ( .A(img[1288]), .B(n28301), .S(n28605), .O(n12244) );
  MUX2S U16076 ( .A(img[1291]), .B(n27668), .S(n28605), .O(n12241) );
  MUX2S U16077 ( .A(img[136]), .B(n28309), .S(n29306), .O(n13396) );
  MUX2S U16078 ( .A(img[139]), .B(n27676), .S(n29306), .O(n13391) );
  MUX2S U16079 ( .A(img[141]), .B(n26557), .S(n29306), .O(n13393) );
  MUX2S U16080 ( .A(img[309]), .B(n26464), .S(n28632), .O(n13225) );
  MUX2S U16081 ( .A(img[533]), .B(n26203), .S(n29021), .O(n13001) );
  MUX2S U16082 ( .A(img[405]), .B(n26243), .S(n29081), .O(n13127) );
  MUX2S U16083 ( .A(img[917]), .B(n26231), .S(n29061), .O(n12615) );
  MUX2S U16084 ( .A(img[789]), .B(n26258), .S(n29102), .O(n12745) );
  MUX2S U16085 ( .A(img[661]), .B(n26262), .S(n29109), .O(n12871) );
  MUX2S U16086 ( .A(img[373]), .B(n26563), .S(n29315), .O(n13161) );
  MUX2S U16087 ( .A(img[293]), .B(n26623), .S(n29361), .O(n13241) );
  MUX2S U16088 ( .A(img[285]), .B(n26077), .S(n29179), .O(n13247) );
  MUX2S U16089 ( .A(img[1165]), .B(n26492), .S(n28590), .O(n12369) );
  MUX2S U16090 ( .A(img[909]), .B(n26553), .S(n29300), .O(n12625) );
  MUX2S U16091 ( .A(img[781]), .B(n26565), .S(n29324), .O(n12751) );
  MUX2S U16092 ( .A(img[653]), .B(n26570), .S(n29331), .O(n12881) );
  MUX2S U16093 ( .A(img[525]), .B(n26549), .S(n29289), .O(n13007) );
  MUX2S U16094 ( .A(img[1725]), .B(n26129), .S(n28948), .O(n11809) );
  MUX2S U16095 ( .A(img[1597]), .B(n26149), .S(n28976), .O(n11935) );
  MUX2S U16096 ( .A(img[21]), .B(n26207), .S(n29027), .O(n13513) );
  MUX2S U16097 ( .A(img[277]), .B(n26239), .S(n29074), .O(n13257) );
  MUX2S U16098 ( .A(img[1461]), .B(n26531), .S(n28652), .O(n12071) );
  MUX2S U16099 ( .A(img[1205]), .B(n26497), .S(n28598), .O(n12327) );
  MUX2S U16100 ( .A(img[1925]), .B(n26186), .S(n29007), .O(n11607) );
  MUX2S U16101 ( .A(img[1797]), .B(n26113), .S(n28906), .O(n11737) );
  MUX2S U16102 ( .A(img[1669]), .B(n26134), .S(n28936), .O(n11863) );
  MUX2S U16103 ( .A(img[1541]), .B(n26155), .S(n28965), .O(n11993) );
  MUX2S U16104 ( .A(img[773]), .B(n26600), .S(n29423), .O(n12761) );
  MUX2S U16105 ( .A(img[645]), .B(n26605), .S(n29430), .O(n12887) );
  MUX2S U16106 ( .A(img[261]), .B(n26578), .S(n29409), .O(n13273) );
  MUX2S U16107 ( .A(img[1173]), .B(n26217), .S(n29040), .O(n12359) );
  MUX2S U16108 ( .A(img[1021]), .B(n26593), .S(n29399), .O(n12513) );
  MUX2S U16109 ( .A(img[973]), .B(n26516), .S(n28623), .O(n12561) );
  MUX2S U16110 ( .A(img[1053]), .B(n26176), .S(n29192), .O(n12479) );
  MUX2S U16111 ( .A(img[77]), .B(n26489), .S(n28587), .O(n13455) );
  MUX2S U16112 ( .A(n26545), .B(img[13]), .S(n29295), .O(n13519) );
  MUX2S U16113 ( .A(n26522), .B(img[437]), .S(n28638), .O(n13095) );
  MUX2S U16114 ( .A(n26635), .B(img[677]), .S(n29380), .O(n12855) );
  MUX2S U16115 ( .A(n26587), .B(img[5]), .S(n29389), .O(n13527) );
  MUX2S U16116 ( .A(n26245), .B(img[1453]), .S(n29087), .O(n12081) );
  MUX2S U16117 ( .A(n26633), .B(img[861]), .S(n29371), .O(n12671) );
  MUX2S U16118 ( .A(n26219), .B(img[1325]), .S(n29047), .O(n12207) );
  MUX2S U16119 ( .A(n26537), .B(img[821]), .S(n28659), .O(n12713) );
  MUX2S U16120 ( .A(n26595), .B(img[389]), .S(n29416), .O(n13143) );
  MUX2S U16121 ( .A(n26118), .B(img[1829]), .S(n28892), .O(n11705) );
  MUX2S U16122 ( .A(img[1160]), .B(n28290), .S(n28590), .O(n12372) );
  MUX2S U16123 ( .A(img[520]), .B(n28276), .S(n29289), .O(n13012) );
  MUX2S U16124 ( .A(img[1338]), .B(n25719), .S(n28835), .O(n12194) );
  MUX2S U16125 ( .A(img[1466]), .B(n25742), .S(n28875), .O(n12062) );
  MUX2S U16126 ( .A(img[1200]), .B(n28282), .S(n28598), .O(n12332) );
  MUX2S U16127 ( .A(img[1922]), .B(n25710), .S(n29007), .O(n11610) );
  MUX2S U16128 ( .A(img[1794]), .B(n25776), .S(n28906), .O(n11734) );
  MUX2S U16129 ( .A(img[642]), .B(n25757), .S(n29430), .O(n12890) );
  MUX2S U16130 ( .A(img[258]), .B(n25733), .S(n29409), .O(n13270) );
  MUX2S U16131 ( .A(img[1818]), .B(n25766), .S(n28899), .O(n11714) );
  MUX2S U16132 ( .A(n28280), .B(img[8]), .S(n29295), .O(n13524) );
  MUX2S U16133 ( .A(n25715), .B(img[514]), .S(n29383), .O(n13014) );
  MUX2S U16134 ( .A(n25761), .B(img[1826]), .S(n28892), .O(n11702) );
  MUX2S U16135 ( .A(img[1163]), .B(n27658), .S(n28590), .O(n12367) );
  MUX2S U16136 ( .A(img[523]), .B(n27644), .S(n29289), .O(n13009) );
  MUX2S U16137 ( .A(img[1595]), .B(n27603), .S(n28976), .O(n11937) );
  MUX2S U16138 ( .A(img[1083]), .B(n27614), .S(n28990), .O(n12449) );
  MUX2S U16139 ( .A(img[1667]), .B(n27577), .S(n28936), .O(n11865) );
  MUX2S U16140 ( .A(img[1539]), .B(n27598), .S(n28965), .O(n11991) );
  MUX2S U16141 ( .A(n27648), .B(img[11]), .S(n29295), .O(n13521) );
  MUX2S U16142 ( .A(img[1007]), .B(n24483), .S(n29064), .O(n12531) );
  MUX2S U16143 ( .A(img[974]), .B(n25191), .S(n28623), .O(n12562) );
  MUX2S U16144 ( .A(img[317]), .B(n26391), .S(n28854), .O(n13215) );
  MUX2S U16145 ( .A(img[1085]), .B(n26419), .S(n28990), .O(n12447) );
  MUX2S U16146 ( .A(img[957]), .B(n26387), .S(n28842), .O(n12577) );
  MUX2S U16147 ( .A(img[1413]), .B(n26399), .S(n28864), .O(n12119) );
  MUX2S U16148 ( .A(img[1285]), .B(n26375), .S(n28824), .O(n12249) );
  MUX2S U16149 ( .A(img[1157]), .B(n26363), .S(n28810), .O(n12375) );
  MUX2S U16150 ( .A(n26409), .B(img[829]), .S(n28883), .O(n12703) );
  MUX2S U16151 ( .A(img[2044]), .B(n29012), .S(n29011), .O(n11488) );
  MUX2S U16152 ( .A(img[1516]), .B(n29100), .S(n29099), .O(n12016) );
  ND2S U16153 ( .I1(n13820), .I2(img[1492]), .O(n29097) );
  MUX2S U16154 ( .A(img[1532]), .B(n28869), .S(n28868), .O(n12000) );
  MUX2S U16155 ( .A(img[1524]), .B(n28650), .S(n28649), .O(n12008) );
  ND2S U16156 ( .I1(n13820), .I2(img[1484]), .O(n28647) );
  MUX2S U16157 ( .A(img[1500]), .B(n29253), .S(n29252), .O(n12032) );
  ND2S U16158 ( .I1(n13820), .I2(img[1508]), .O(n29250) );
  MUX2S U16159 ( .A(img[1884]), .B(n28897), .S(n28896), .O(n11648) );
  MUX2S U16160 ( .A(img[1756]), .B(n28927), .S(n28926), .O(n11776) );
  MUX2S U16161 ( .A(img[1628]), .B(n28956), .S(n28955), .O(n11904) );
  ND2S U16162 ( .I1(n13820), .I2(img[1228]), .O(n28593) );
  ND2S U16163 ( .I1(n13819), .I2(img[1220]), .O(n28812) );
  ND2S U16164 ( .I1(n13820), .I2(img[1900]), .O(n28674) );
  ND2S U16165 ( .I1(n13819), .I2(img[1380]), .O(n29235) );
  ND2S U16166 ( .I1(n13820), .I2(img[1396]), .O(n28615) );
  ND2S U16167 ( .I1(n13820), .I2(img[1244]), .O(n29216) );
  ND2S U16168 ( .I1(n13820), .I2(img[2036]), .O(n28794) );
  ND2S U16169 ( .I1(n13819), .I2(img[1908]), .O(n28696) );
  ND2S U16170 ( .I1(n13905), .I2(img[1140]), .O(n28766) );
  ND2S U16171 ( .I1(n13819), .I2(img[1260]), .O(n29035) );
  MUX2S U16172 ( .A(img[2046]), .B(n24943), .S(n29011), .O(n11486) );
  MUX2S U16173 ( .A(img[2041]), .B(n26821), .S(n29011), .O(n11491) );
  MUX2S U16174 ( .A(img[904]), .B(n28305), .S(n29300), .O(n12628) );
  MUX2S U16175 ( .A(img[907]), .B(n27672), .S(n29300), .O(n12623) );
  MUX2S U16176 ( .A(img[651]), .B(n27705), .S(n29331), .O(n12879) );
  MUX2S U16177 ( .A(img[1527]), .B(n23988), .S(n28649), .O(n12005) );
  ND2S U16178 ( .I1(n29258), .I2(img[1487]), .O(n23985) );
  MUX2S U16179 ( .A(img[1503]), .B(n24197), .S(n29252), .O(n12035) );
  ND2S U16180 ( .I1(n13819), .I2(img[1511]), .O(n24194) );
  MUX2S U16181 ( .A(img[1887]), .B(n24245), .S(n28896), .O(n11645) );
  ND2S U16182 ( .I1(n13820), .I2(img[1895]), .O(n24242) );
  MUX2S U16183 ( .A(img[1759]), .B(n24272), .S(n28926), .O(n11779) );
  ND2S U16184 ( .I1(n29124), .I2(img[1767]), .O(n24269) );
  MUX2S U16185 ( .A(img[1631]), .B(n24299), .S(n28955), .O(n11901) );
  ND2S U16186 ( .I1(n13904), .I2(img[1231]), .O(n23920) );
  ND2S U16187 ( .I1(n13819), .I2(img[1223]), .O(n24363) );
  ND2S U16188 ( .I1(n13905), .I2(img[1255]), .O(n24150) );
  ND2S U16189 ( .I1(n13819), .I2(img[1407]), .O(n24381) );
  ND2S U16190 ( .I1(n13904), .I2(img[1375]), .O(n24166) );
  ND2S U16191 ( .I1(n29124), .I2(img[1655]), .O(n24093) );
  ND2S U16192 ( .I1(n13819), .I2(img[1391]), .O(n24471) );
  ND2S U16193 ( .I1(n13819), .I2(img[1399]), .O(n23947) );
  ND2S U16194 ( .I1(n13905), .I2(img[1903]), .O(n24017) );
  ND2S U16195 ( .I1(n29124), .I2(img[1791]), .O(n24256) );
  ND2S U16196 ( .I1(n13819), .I2(img[1095]), .O(n24435) );
  ND2S U16197 ( .I1(n13904), .I2(img[1111]), .O(n24539) );
  ND2S U16198 ( .I1(n13904), .I2(img[1143]), .O(n24107) );
  ND2S U16199 ( .I1(n13819), .I2(img[1783]), .O(n24069) );
  MUX2S U16200 ( .A(img[1521]), .B(n27142), .S(n28649), .O(n12011) );
  ND2S U16201 ( .I1(n13902), .I2(img[1481]), .O(n27140) );
  MUX2S U16202 ( .A(img[1526]), .B(n25005), .S(n28649), .O(n12006) );
  ND2S U16203 ( .I1(n13901), .I2(img[1486]), .O(n25003) );
  MUX2S U16204 ( .A(img[2009]), .B(n26808), .S(n28997), .O(n11517) );
  MUX2S U16205 ( .A(img[2014]), .B(n24933), .S(n28997), .O(n11522) );
  ND2S U16206 ( .I1(n13900), .I2(img[2022]), .O(n24931) );
  MUX2S U16207 ( .A(img[1529]), .B(n26723), .S(n28868), .O(n11997) );
  MUX2S U16208 ( .A(img[1497]), .B(n26875), .S(n29252), .O(n12029) );
  MUX2S U16209 ( .A(img[1502]), .B(n25154), .S(n29252), .O(n12034) );
  ND2S U16210 ( .I1(n13819), .I2(img[1510]), .O(n25152) );
  MUX2S U16211 ( .A(img[1758]), .B(n24882), .S(n28926), .O(n11778) );
  MUX2S U16212 ( .A(img[1630]), .B(n24903), .S(n28955), .O(n11902) );
  ND2S U16213 ( .I1(n13819), .I2(img[1638]), .O(n24901) );
  ND2S U16214 ( .I1(n13819), .I2(img[1353]), .O(n27118) );
  ND2S U16215 ( .I1(n29124), .I2(img[1217]), .O(n26684) );
  ND2S U16216 ( .I1(n13770), .I2(img[2030]), .O(n25088) );
  ND2S U16217 ( .I1(n29124), .I2(img[1918]), .O(n24875) );
  ND2S U16218 ( .I1(n13903), .I2(img[1657]), .O(n26786) );
  ND2S U16219 ( .I1(n13903), .I2(img[1662]), .O(n24916) );
  ND2S U16220 ( .I1(n13903), .I2(img[1350]), .O(n24814) );
  ND2S U16221 ( .I1(n13904), .I2(img[1129]), .O(n27062) );
  ND2S U16222 ( .I1(n13903), .I2(img[1390]), .O(n25286) );
  ND2S U16223 ( .I1(n13903), .I2(img[1910]), .O(n25027) );
  ND2S U16224 ( .I1(n13770), .I2(img[2025]), .O(n27084) );
  ND2S U16225 ( .I1(n13903), .I2(img[1150]), .O(n24926) );
  ND2S U16226 ( .I1(n13819), .I2(img[1110]), .O(n25304) );
  ND2S U16227 ( .I1(n13770), .I2(img[1121]), .O(n26892) );
  ND2S U16228 ( .I1(n13902), .I2(img[1126]), .O(n25172) );
  ND2S U16229 ( .I1(n29124), .I2(img[1137]), .O(n27149) );
  ND2S U16230 ( .I1(n13820), .I2(img[1142]), .O(n25078) );
  ND2S U16231 ( .I1(n13903), .I2(img[1905]), .O(n26996) );
  ND2S U16232 ( .I1(n13904), .I2(img[1641]), .O(n27052) );
  ND2S U16233 ( .I1(n13905), .I2(img[1646]), .O(n25057) );
  ND2S U16234 ( .I1(n13903), .I2(img[1777]), .O(n27016) );
  MUX2S U16235 ( .A(img[1507]), .B(n27804), .S(n29261), .O(n12025) );
  ND2S U16236 ( .I1(n13819), .I2(img[1499]), .O(n27802) );
  MUX2S U16237 ( .A(img[1883]), .B(n27550), .S(n28896), .O(n11649) );
  MUX2S U16238 ( .A(img[1755]), .B(n27570), .S(n28926), .O(n11775) );
  ND2S U16239 ( .I1(n13903), .I2(img[1763]), .O(n27568) );
  ND2S U16240 ( .I1(n13903), .I2(img[1915]), .O(n27563) );
  ND2S U16241 ( .I1(n29124), .I2(img[1787]), .O(n27583) );
  ND2S U16242 ( .I1(n13903), .I2(img[1123]), .O(n27762) );
  ND2S U16243 ( .I1(n13903), .I2(img[1131]), .O(n27419) );
  ND2S U16244 ( .I1(n13903), .I2(img[1139]), .O(n27708) );
  ND2S U16245 ( .I1(n13903), .I2(img[1371]), .O(n27784) );
  ND2S U16246 ( .I1(n29258), .I2(img[1243]), .O(n27774) );
  ND2S U16247 ( .I1(n13903), .I2(img[1347]), .O(n27501) );
  ND2S U16248 ( .I1(n13903), .I2(img[1219]), .O(n27491) );
  ND2S U16249 ( .I1(n13903), .I2(img[2035]), .O(n27429) );
  ND2S U16250 ( .I1(n13819), .I2(img[1771]), .O(n27389) );
  ND2S U16251 ( .I1(n13903), .I2(img[1651]), .O(n27399) );
  ND2S U16252 ( .I1(n13903), .I2(img[1387]), .O(n27310) );
  ND2S U16253 ( .I1(n13819), .I2(img[1395]), .O(n27661) );
  ND2S U16254 ( .I1(n13903), .I2(img[1531]), .O(n27533) );
  ND2S U16255 ( .I1(n13903), .I2(img[1259]), .O(n27300) );
  MUX2S U16256 ( .A(img[2040]), .B(n28072), .S(n29011), .O(n11492) );
  MUX2S U16257 ( .A(img[1520]), .B(n28326), .S(n28649), .O(n12012) );
  ND2S U16258 ( .I1(n13819), .I2(img[1480]), .O(n28324) );
  MUX2S U16259 ( .A(img[1498]), .B(n25919), .S(n29252), .O(n12030) );
  ND2S U16260 ( .I1(n13819), .I2(img[1506]), .O(n25917) );
  MUX2S U16261 ( .A(img[2010]), .B(n25698), .S(n28997), .O(n11518) );
  MUX2S U16262 ( .A(img[2008]), .B(n28061), .S(n28997), .O(n11524) );
  ND2S U16263 ( .I1(n13904), .I2(img[2016]), .O(n28059) );
  MUX2S U16264 ( .A(img[1528]), .B(n27956), .S(n28868), .O(n12004) );
  ND2S U16265 ( .I1(n13819), .I2(img[1472]), .O(n27954) );
  MUX2S U16266 ( .A(img[1530]), .B(n25750), .S(n28868), .O(n11998) );
  ND2S U16267 ( .I1(n13904), .I2(img[1474]), .O(n25748) );
  MUX2S U16268 ( .A(img[1512]), .B(n28170), .S(n29099), .O(n12020) );
  ND2S U16269 ( .I1(n13819), .I2(img[1488]), .O(n28168) );
  MUX2S U16270 ( .A(img[1496]), .B(n28404), .S(n29252), .O(n12036) );
  ND2S U16271 ( .I1(n13819), .I2(img[1504]), .O(n28402) );
  MUX2S U16272 ( .A(img[1752]), .B(n28009), .S(n28926), .O(n11780) );
  MUX2S U16273 ( .A(img[1624]), .B(n28029), .S(n28955), .O(n11908) );
  ND2S U16274 ( .I1(n13904), .I2(img[1240]), .O(n28360) );
  ND2S U16275 ( .I1(n13904), .I2(img[2026]), .O(n25558) );
  ND2S U16276 ( .I1(n13819), .I2(img[2034]), .O(n25568) );
  ND2S U16277 ( .I1(n13904), .I2(img[1370]), .O(n25889) );
  ND2S U16278 ( .I1(n13819), .I2(img[1904]), .O(n28183) );
  ND2S U16279 ( .I1(n13904), .I2(img[1344]), .O(n27969) );
  ND2S U16280 ( .I1(n13819), .I2(img[1346]), .O(n25725) );
  ND2S U16281 ( .I1(n13904), .I2(img[1138]), .O(n25548) );
  ND2S U16282 ( .I1(n13819), .I2(img[1362]), .O(n25598) );
  ND2S U16283 ( .I1(n13904), .I2(img[1640]), .O(n28234) );
  ND2S U16284 ( .I1(n13819), .I2(img[1648]), .O(n28224) );
  ND2S U16285 ( .I1(n13819), .I2(img[1384]), .O(n28136) );
  ND2S U16286 ( .I1(n13900), .I2(img[1906]), .O(n25498) );
  ND2S U16287 ( .I1(n13900), .I2(img[1234]), .O(n25586) );
  ND2S U16288 ( .I1(n13904), .I2(img[1784]), .O(n28022) );
  ND2S U16289 ( .I1(n13904), .I2(img[1106]), .O(n25643) );
  ND2S U16290 ( .I1(n13900), .I2(img[1122]), .O(n25936) );
  ND2S U16291 ( .I1(n13900), .I2(img[1256]), .O(n28125) );
  ND2S U16292 ( .I1(n13904), .I2(img[2042]), .O(n25706) );
  ND2S U16293 ( .I1(n13904), .I2(img[1522]), .O(n25469) );
  MUX2S U16294 ( .A(img[356]), .B(n29183), .S(n29182), .O(n13176) );
  MUX2S U16295 ( .A(img[340]), .B(n29158), .S(n29157), .O(n13192) );
  MUX2S U16296 ( .A(img[1517]), .B(n26251), .S(n29099), .O(n12017) );
  MUX2S U16297 ( .A(img[1501]), .B(n26088), .S(n29252), .O(n12033) );
  MUX2S U16298 ( .A(n29186), .B(img[1060]), .S(n29185), .O(n12472) );
  MUX2S U16299 ( .A(img[1629]), .B(n26163), .S(n28955), .O(n11903) );
  ND2S U16300 ( .I1(n13900), .I2(img[1637]), .O(n26161) );
  MUX2S U16301 ( .A(img[2013]), .B(n26194), .S(n28997), .O(n11521) );
  ND2S U16302 ( .I1(n13900), .I2(img[2021]), .O(n26192) );
  MUX2S U16303 ( .A(img[1525]), .B(n26529), .S(n28649), .O(n12007) );
  MUX2S U16304 ( .A(n29167), .B(img[812]), .S(n29166), .O(n12720) );
  MUX2S U16305 ( .A(img[1757]), .B(n26142), .S(n28926), .O(n11777) );
  ND2S U16306 ( .I1(n13904), .I2(img[1909]), .O(n26265) );
  ND2S U16307 ( .I1(n13900), .I2(img[1245]), .O(n26055) );
  ND2S U16308 ( .I1(n13904), .I2(img[1357]), .O(n26505) );
  ND2S U16309 ( .I1(n13900), .I2(img[1901]), .O(n26275) );
  ND2S U16310 ( .I1(n13900), .I2(img[1381]), .O(n26060) );
  ND2S U16311 ( .I1(n13904), .I2(img[1645]), .O(n26315) );
  ND2S U16312 ( .I1(n13900), .I2(img[1653]), .O(n26305) );
  ND2S U16313 ( .I1(n13904), .I2(img[1773]), .O(n26295) );
  ND2S U16314 ( .I1(n13900), .I2(img[1093]), .O(n26415) );
  ND2S U16315 ( .I1(n13904), .I2(img[1125]), .O(n26172) );
  ND2S U16316 ( .I1(n13900), .I2(img[1261]), .O(n26210) );
  ND2S U16317 ( .I1(n13904), .I2(img[1781]), .O(n26285) );
  MUX2S U16318 ( .A(n27035), .B(img[1585]), .S(n28750), .O(n11941) );
  MUX2S U16319 ( .A(n27056), .B(img[1041]), .S(n29122), .O(n12491) );
  MUX2S U16320 ( .A(img[535]), .B(n24450), .S(n29021), .O(n13003) );
  MUX2S U16321 ( .A(img[23]), .B(n24454), .S(n29027), .O(n13515) );
  MUX2S U16322 ( .A(img[279]), .B(n24496), .S(n29074), .O(n13259) );
  MUX2S U16323 ( .A(img[1175]), .B(n24467), .S(n29040), .O(n12357) );
  MUX2S U16324 ( .A(img[1431]), .B(n24521), .S(n29094), .O(n12101) );
  MUX2S U16325 ( .A(img[1199]), .B(n24456), .S(n29033), .O(n12339) );
  MUX2S U16326 ( .A(img[334]), .B(n25199), .S(n28635), .O(n13198) );
  MUX2S U16327 ( .A(img[54]), .B(n25185), .S(n28584), .O(n13479) );
  MUX2S U16328 ( .A(img[1054]), .B(n25179), .S(n29192), .O(n12478) );
  MUX2S U16329 ( .A(img[94]), .B(n25220), .S(n29339), .O(n13438) );
  MUX2S U16330 ( .A(img[113]), .B(n27109), .S(n29536), .O(n13413) );
  MUX2S U16331 ( .A(img[371]), .B(n27678), .S(n29315), .O(n13159) );
  MUX2S U16332 ( .A(img[51]), .B(n27717), .S(n28584), .O(n13481) );
  MUX2S U16333 ( .A(n25832), .B(img[2]), .S(n29389), .O(n13530) );
  MUX2S U16334 ( .A(n25801), .B(img[1570]), .S(n28951), .O(n11958) );
  MUX2S U16335 ( .A(n28339), .B(img[1072]), .S(n28764), .O(n12460) );
  MUX2S U16336 ( .A(img[2012]), .B(n28998), .S(n28997), .O(n11520) );
  ND2S U16337 ( .I1(n13901), .I2(img[2020]), .O(n28995) );
  MUX2S U16338 ( .A(img[368]), .B(n28311), .S(n29315), .O(n13164) );
  ND2S U16339 ( .I1(n13901), .I2(img[1660]), .O(n28971) );
  ND2S U16340 ( .I1(n13904), .I2(img[1116]), .O(n29195) );
  ND2S U16341 ( .I1(n13904), .I2(img[1348]), .O(n28826) );
  MUX2S U16342 ( .A(img[1666]), .B(n25796), .S(n28936), .O(n11866) );
  MUX2S U16343 ( .A(img[1538]), .B(n25817), .S(n28965), .O(n11990) );
  ND2S U16344 ( .I1(n13901), .I2(img[1788]), .O(n28943) );
  MUX2S U16345 ( .A(img[1456]), .B(n28320), .S(n28652), .O(n12076) );
  MUX2S U16346 ( .A(img[1562]), .B(n25806), .S(n28958), .O(n11970) );
  MUX2S U16347 ( .A(img[1722]), .B(n25791), .S(n28948), .O(n11806) );
  MUX2S U16348 ( .A(img[1594]), .B(n25812), .S(n28976), .O(n11938) );
  MUX2S U16349 ( .A(img[1026]), .B(n25827), .S(n28979), .O(n12502) );
  MUX2S U16350 ( .A(img[1082]), .B(n25822), .S(n28990), .O(n12450) );
  MUX2S U16351 ( .A(img[1690]), .B(n25786), .S(n28929), .O(n11838) );
  MUX2S U16352 ( .A(img[32]), .B(n28355), .S(n29342), .O(n13500) );
  MUX2S U16353 ( .A(img[898]), .B(n25836), .S(n29395), .O(n12634) );
  MUX2S U16354 ( .A(img[2015]), .B(n24342), .S(n28997), .O(n11523) );
  ND2S U16355 ( .I1(n13904), .I2(img[2023]), .O(n24338) );
  ND2S U16356 ( .I1(n13901), .I2(img[1127]), .O(n24310) );
  ND2S U16357 ( .I1(n13901), .I2(img[1647]), .O(n24074) );
  MUX2S U16358 ( .A(img[1753]), .B(n26758), .S(n28926), .O(n11773) );
  ND2S U16359 ( .I1(n13901), .I2(img[1761]), .O(n26756) );
  MUX2S U16360 ( .A(img[1625]), .B(n26778), .S(n28955), .O(n11907) );
  ND2S U16361 ( .I1(n13901), .I2(img[1633]), .O(n26776) );
  ND2S U16362 ( .I1(n13904), .I2(img[1233]), .O(n26940) );
  ND2S U16363 ( .I1(n13904), .I2(img[1361]), .O(n26950) );
  ND2S U16364 ( .I1(n13904), .I2(img[2033]), .O(n27068) );
  MUX2S U16365 ( .A(img[1886]), .B(n24862), .S(n28896), .O(n11646) );
  ND2S U16366 ( .I1(n13901), .I2(img[1089]), .O(n26799) );
  ND2S U16367 ( .I1(n13901), .I2(img[1246]), .O(n25119) );
  ND2S U16368 ( .I1(n13901), .I2(img[1382]), .O(n25126) );
  ND2S U16369 ( .I1(n13901), .I2(img[2038]), .O(n25098) );
  ND2S U16370 ( .I1(n13901), .I2(img[1262]), .O(n25325) );
  ND2S U16371 ( .I1(n13904), .I2(img[1534]), .O(n24845) );
  MUX2S U16372 ( .A(img[2047]), .B(n24333), .S(n29011), .O(n13533) );
  ND3S U16373 ( .I1(n24340), .I2(n24329), .I3(n24328), .O(n24333) );
  ND3S U16374 ( .I1(n27070), .I2(n26742), .I3(n26741), .O(n26743) );
  MUX2S U16375 ( .A(img[341]), .B(n26450), .S(n29157), .O(n13193) );
  MUX2S U16376 ( .A(n26456), .B(img[813]), .S(n29166), .O(n12719) );
  MUX2S U16377 ( .A(n26984), .B(img[1489]), .S(n29091), .O(n12043) );
  ND3S U16378 ( .I1(n27170), .I2(n26983), .I3(n26982), .O(n26984) );
  MUX2S U16379 ( .A(n25299), .B(img[1494]), .S(n29091), .O(n12038) );
  ND3S U16380 ( .I1(n25298), .I2(n25297), .I3(n25296), .O(n25299) );
  ND2S U16381 ( .I1(n13901), .I2(img[1518]), .O(n25296) );
  MUX2S U16382 ( .A(n24512), .B(img[1495]), .S(n29091), .O(n12037) );
  ND3S U16383 ( .I1(n24581), .I2(n24507), .I3(n24506), .O(n24512) );
  ND2S U16384 ( .I1(n13904), .I2(img[1519]), .O(n24506) );
  ND2S U16385 ( .I1(n13902), .I2(img[1533]), .O(n26405) );
  MUX2S U16386 ( .A(img[1627]), .B(n27591), .S(n28955), .O(n11905) );
  ND2S U16387 ( .I1(n13902), .I2(img[1635]), .O(n27589) );
  MUX2S U16388 ( .A(img[2027]), .B(n27446), .S(n28782), .O(n11503) );
  MUX2S U16389 ( .A(img[2019]), .B(n27630), .S(n29004), .O(n11513) );
  MUX2S U16390 ( .A(img[1739]), .B(n27381), .S(n28726), .O(n11791) );
  ND2S U16391 ( .I1(n13902), .I2(img[1515]), .O(n27337) );
  MUX2S U16392 ( .A(img[1907]), .B(n27364), .S(n28690), .O(n11623) );
  MUX2S U16393 ( .A(img[1483]), .B(n27691), .S(n28656), .O(n12047) );
  ND2S U16394 ( .I1(n13902), .I2(img[1523]), .O(n27689) );
  MUX2S U16395 ( .A(img[1147]), .B(n27612), .S(n28983), .O(n12385) );
  ND2S U16396 ( .I1(n13902), .I2(img[1091]), .O(n27610) );
  MUX2S U16397 ( .A(n25740), .B(img[506]), .S(n29420), .O(n13022) );
  MUX2S U16398 ( .A(n26713), .B(img[505]), .S(n29420), .O(n13021) );
  MUX2S U16399 ( .A(n25250), .B(img[510]), .S(n29420), .O(n13026) );
  MUX2S U16400 ( .A(n28102), .B(img[504]), .S(n29420), .O(n13028) );
  MUX2S U16401 ( .A(n24742), .B(img[511]), .S(n29420), .O(n13027) );
  ND2S U16402 ( .I1(n13904), .I2(img[2037]), .O(n26336) );
  ND2S U16403 ( .I1(n13902), .I2(img[1141]), .O(n26475) );
  ND2S U16404 ( .I1(n13902), .I2(img[1917]), .O(n26109) );
  ND2S U16405 ( .I1(n13904), .I2(img[1405]), .O(n26383) );
  MUX2S U16406 ( .A(n26989), .B(img[849]), .S(n29170), .O(n12677) );
  MUX2S U16407 ( .A(n25755), .B(img[890]), .S(n29427), .O(n12642) );
  MUX2S U16408 ( .A(n26880), .B(img[857]), .S(n29371), .O(n12675) );
  MUX2S U16409 ( .A(n25681), .B(img[874]), .S(n29106), .O(n12658) );
  MUX2S U16410 ( .A(n24630), .B(img[863]), .S(n29371), .O(n12669) );
  MUX2S U16411 ( .A(n27255), .B(img[873]), .S(n29106), .O(n12659) );
  MUX2S U16412 ( .A(n28489), .B(img[840]), .S(n28663), .O(n12692) );
  MUX2S U16413 ( .A(n25924), .B(img[858]), .S(n29371), .O(n12674) );
  MUX2S U16414 ( .A(n24208), .B(img[871]), .S(n29230), .O(n12667) );
  MUX2S U16415 ( .A(n27101), .B(img[881]), .S(n29328), .O(n12645) );
  MUX2S U16416 ( .A(n27538), .B(img[827]), .S(n28883), .O(n12705) );
  MUX2S U16417 ( .A(n28522), .B(img[864]), .S(n29230), .O(n12668) );
  MUX2S U16418 ( .A(n24573), .B(img[855]), .S(n29170), .O(n12683) );
  MUX2S U16419 ( .A(n23999), .B(img[847]), .S(n28663), .O(n12685) );
  MUX2S U16420 ( .A(n24751), .B(img[895]), .S(n29427), .O(n12637) );
  MUX2S U16421 ( .A(n28409), .B(img[856]), .S(n29371), .O(n12676) );
  MUX2S U16422 ( .A(n25162), .B(img[870]), .S(n29230), .O(n12666) );
  MUX2S U16423 ( .A(n25010), .B(img[886]), .S(n29328), .O(n12650) );
  MUX2S U16424 ( .A(n24679), .B(img[887]), .S(n29328), .O(n12651) );
  MUX2S U16425 ( .A(n26003), .B(img[826]), .S(n28883), .O(n12706) );
  MUX2S U16426 ( .A(n28108), .B(img[888]), .S(n29427), .O(n12644) );
  MUX2S U16427 ( .A(n25636), .B(img[850]), .S(n29170), .O(n12678) );
  MUX2S U16428 ( .A(n28175), .B(img[872]), .S(n29106), .O(n12660) );
  MUX2S U16429 ( .A(n28455), .B(img[848]), .S(n29170), .O(n12684) );
  MUX2S U16430 ( .A(n27224), .B(img[825]), .S(n28883), .O(n12707) );
  MUX2S U16431 ( .A(n25386), .B(img[878]), .S(n29106), .O(n12654) );
  MUX2S U16432 ( .A(n28331), .B(img[880]), .S(n29328), .O(n12652) );
  MUX2S U16433 ( .A(n25350), .B(img[854]), .S(n29170), .O(n12682) );
  MUX2S U16434 ( .A(n27850), .B(img[891]), .S(n29427), .O(n12641) );
  MUX2S U16435 ( .A(n26923), .B(img[865]), .S(n29230), .O(n12661) );
  MUX2S U16436 ( .A(n25864), .B(img[842]), .S(n28663), .O(n12690) );
  MUX2S U16437 ( .A(n25276), .B(img[894]), .S(n29427), .O(n12638) );
  MUX2S U16438 ( .A(n24418), .B(img[831]), .S(n28883), .O(n12701) );
  MUX2S U16439 ( .A(n25241), .B(img[862]), .S(n29371), .O(n12670) );
  MUX2S U16440 ( .A(n24853), .B(img[838]), .S(n28879), .O(n12698) );
  MUX2S U16441 ( .A(n24525), .B(img[879]), .S(n29106), .O(n12653) );
  MUX2S U16442 ( .A(n25208), .B(img[846]), .S(n28663), .O(n12686) );
  MUX2S U16443 ( .A(n27699), .B(img[883]), .S(n29328), .O(n12647) );
  MUX2S U16444 ( .A(n25479), .B(img[882]), .S(n29328), .O(n12646) );
  MUX2S U16445 ( .A(n27997), .B(img[824]), .S(n28883), .O(n12708) );
  ND2S U16446 ( .I1(n23121), .I2(n23120), .O(n23126) );
  ND2S U16447 ( .I1(n23133), .I2(n23132), .O(n23136) );
  ND2S U16448 ( .I1(n23359), .I2(n23364), .O(n23367) );
  ND2S U16449 ( .I1(n23386), .I2(n23385), .O(n23388) );
  ND2S U16450 ( .I1(n23397), .I2(n23396), .O(n23398) );
  XOR3S U16451 ( .I1(n21802), .I2(n21801), .I3(mult_x_431_n11), .O(PE_N56) );
  ND2S U16452 ( .I1(n22402), .I2(n22401), .O(mult_x_433_n8) );
  XOR3S U16453 ( .I1(n22402), .I2(n22401), .I3(mult_x_433_n9), .O(PE_N90) );
  XOR3S U16454 ( .I1(n22404), .I2(n22403), .I3(mult_x_433_n14), .O(PE_N88) );
  ND2S U16455 ( .I1(n22610), .I2(n22609), .O(n22612) );
  ND2S U16456 ( .I1(n22615), .I2(n22614), .O(n22618) );
  ND2S U16457 ( .I1(n22626), .I2(n22625), .O(n22627) );
  ND2S U16458 ( .I1(n22000), .I2(n21999), .O(n22002) );
  ND2S U16459 ( .I1(n22252), .I2(n22251), .O(n22254) );
  ND2S U16460 ( .I1(n30026), .I2(n23691), .O(n14011) );
  MXL2HS U16461 ( .A(n21548), .B(n21547), .S(gray_avg[7]), .OB(gray_avg[6]) );
  OR2S U16462 ( .I1(n13926), .I2(n21546), .O(n21547) );
  MXL2HS U16463 ( .A(n21576), .B(n21575), .S(gray_avg[5]), .OB(gray_avg[4]) );
  OR2S U16464 ( .I1(n13918), .I2(n21574), .O(n21575) );
  MXL2HS U16465 ( .A(n23443), .B(n23442), .S(gray_avg[3]), .OB(gray_avg[2]) );
  OR2S U16466 ( .I1(n13922), .I2(n23441), .O(n23442) );
  MUX2S U16467 ( .A(n13919), .B(n23467), .S(gray_avg[1]), .O(gray_avg[0]) );
  MUX2S U16468 ( .A(n29957), .B(rgb_value[6]), .S(n29956), .O(gray_max[6]) );
  MUX2S U16469 ( .A(n29954), .B(rgb_value[5]), .S(n29956), .O(gray_max[5]) );
  MUX2S U16470 ( .A(n29952), .B(rgb_value[4]), .S(n29956), .O(gray_max[4]) );
  MUX2S U16471 ( .A(n29950), .B(rgb_value[3]), .S(n29956), .O(gray_max[3]) );
  MUX2S U16472 ( .A(n29948), .B(rgb_value[2]), .S(n29956), .O(gray_max[2]) );
  MUX2S U16473 ( .A(n29946), .B(rgb_value[1]), .S(n29956), .O(gray_max[1]) );
  MUX2S U16474 ( .A(n29944), .B(rgb_value[0]), .S(n29956), .O(gray_max[0]) );
  INV3 U16475 ( .I(n18297), .O(n15751) );
  NR2 U16476 ( .I1(n14033), .I2(n23624), .O(n16001) );
  ND2 U16477 ( .I1(n14056), .I2(n14045), .O(n16009) );
  INV2 U16478 ( .I(n14077), .O(n15809) );
  BUF1 U16479 ( .I(n13886), .O(n19252) );
  INV4 U16480 ( .I(n15277), .O(n15752) );
  BUF3 U16481 ( .I(n14111), .O(n15653) );
  BUF2 U16482 ( .I(n16001), .O(n14266) );
  INV1S U16483 ( .I(n16364), .O(n16375) );
  INV3 U16484 ( .I(n14299), .O(n17088) );
  INV2 U16485 ( .I(n13929), .O(n20263) );
  INV2 U16486 ( .I(n17658), .O(n17928) );
  INV3 U16487 ( .I(n13927), .O(n17938) );
  BUF1CK U16488 ( .I(n14111), .O(n14112) );
  BUF3 U16489 ( .I(n16364), .O(n14392) );
  BUF2 U16490 ( .I(n16364), .O(n16799) );
  INV2 U16491 ( .I(n13872), .O(n18681) );
  INV2 U16492 ( .I(n17522), .O(n17115) );
  INV2 U16493 ( .I(n16431), .O(n16758) );
  INV1S U16494 ( .I(n18297), .O(n18934) );
  INV2 U16495 ( .I(n17885), .O(n14555) );
  INV1S U16496 ( .I(n14299), .O(n17828) );
  INV2 U16497 ( .I(n16059), .O(n17762) );
  INV1S U16498 ( .I(n16758), .O(n19318) );
  OA112S U16499 ( .C1(n21467), .C2(n29504), .A1(n21466), .B1(n21465), .O(
        n13907) );
  AN2 U16500 ( .I1(n16178), .I2(n16177), .O(n13910) );
  NR2T U16501 ( .I1(n23895), .I2(n14017), .O(n13911) );
  BUF2 U16502 ( .I(n13886), .O(n19641) );
  OA12 U16503 ( .B1(n22942), .B2(n22941), .A1(n22940), .O(n13913) );
  INV2 U16504 ( .I(n21245), .O(n23508) );
  BUF2 U16505 ( .I(n17514), .O(n17617) );
  BUF1CK U16506 ( .I(n19573), .O(n20345) );
  BUF1 U16507 ( .I(n15568), .O(n17730) );
  BUF1S U16508 ( .I(n13800), .O(n17589) );
  BUF1S U16509 ( .I(n13800), .O(n18713) );
  BUF1S U16510 ( .I(n13800), .O(n17612) );
  BUF1S U16511 ( .I(n13800), .O(n18818) );
  BUF1 U16512 ( .I(n19710), .O(n19289) );
  BUF2 U16513 ( .I(n17418), .O(n19914) );
  AOI12HS U16514 ( .B1(n22923), .B2(n22920), .A1(n22919), .O(n13915) );
  AOI12HS U16515 ( .B1(n22923), .B2(n22922), .A1(n22921), .O(n13916) );
  BUF1S U16516 ( .I(n20039), .O(n19955) );
  BUF1S U16517 ( .I(n15561), .O(n19417) );
  BUF1S U16518 ( .I(n15568), .O(n18702) );
  BUF1S U16519 ( .I(n15561), .O(n19349) );
  BUF1S U16520 ( .I(n15561), .O(n17712) );
  BUF1S U16521 ( .I(n20039), .O(n17865) );
  BUF1S U16522 ( .I(n15561), .O(n18838) );
  OAI12HS U16523 ( .B1(n23508), .B2(n19438), .A1(n19058), .O(n19059) );
  BUF1S U16524 ( .I(n15561), .O(n18974) );
  BUF1S U16525 ( .I(n20039), .O(n17767) );
  BUF1S U16526 ( .I(n15561), .O(n18623) );
  BUF1S U16527 ( .I(n15561), .O(n17276) );
  OR2 U16528 ( .I1(i_col[0]), .I2(n14227), .O(n19462) );
  BUF1S U16529 ( .I(n20039), .O(n19295) );
  BUF1S U16530 ( .I(n20039), .O(n19271) );
  BUF1S U16531 ( .I(n15561), .O(n17745) );
  BUF1S U16532 ( .I(n15561), .O(n17840) );
  BUF1S U16533 ( .I(n15561), .O(n19319) );
  INV1S U16534 ( .I(n21669), .O(n22324) );
  INV1S U16535 ( .I(n23770), .O(n29526) );
  BUF1 U16536 ( .I(n28318), .O(n26855) );
  XOR2HS U16537 ( .I1(img_size[3]), .I2(n23954), .O(n23795) );
  ND2S U16538 ( .I1(n21470), .I2(n21430), .O(n21429) );
  OAI222S U16539 ( .A1(n21652), .A2(n21651), .B1(n23770), .B2(n21650), .C1(
        n27893), .C2(n21503), .O(n11261) );
  OAI222S U16540 ( .A1(n21626), .A2(n21651), .B1(n23770), .B2(n21625), .C1(
        n21624), .C2(n21503), .O(n11389) );
  OAI222S U16541 ( .A1(n21609), .A2(n21651), .B1(n23770), .B2(n21608), .C1(
        n21607), .C2(n21503), .O(n11421) );
  INV3 U16542 ( .I(n22060), .O(n17195) );
  AO13 U16543 ( .B1(n22928), .B2(n22927), .B3(n13887), .A1(n22926), .O(n22929)
         );
  OR2P U16544 ( .I1(n22928), .I2(n13910), .O(n18133) );
  INV2 U16545 ( .I(n22928), .O(n14053) );
  NR2 U16546 ( .I1(n15323), .I2(n15322), .O(n15324) );
  NR2 U16547 ( .I1(n15200), .I2(n15199), .O(n15201) );
  NR3 U16548 ( .I1(n15617), .I2(n15616), .I3(n15615), .O(n15624) );
  NR2P U16549 ( .I1(n13844), .I2(n19473), .O(n20366) );
  NR2P U16550 ( .I1(n18134), .I2(n19473), .O(n19601) );
  NR2T U16551 ( .I1(n18132), .I2(n19473), .O(n20363) );
  AOI12HS U16552 ( .B1(n17957), .B2(n20364), .A1(n17956), .O(n17959) );
  AOI12HP U16553 ( .B1(n26039), .B2(n28575), .A1(n26038), .O(n26583) );
  MOAI1 U16554 ( .A1(n20917), .A2(n20916), .B1(n21474), .B2(n21428), .O(n20918) );
  OAI12HS U16555 ( .B1(n28536), .B2(n21607), .A1(n26016), .O(n26039) );
  INV3 U16556 ( .I(n19494), .O(n22922) );
  AN4 U16557 ( .I1(n17129), .I2(n17128), .I3(n17127), .I4(n17126), .O(n17130)
         );
  AOI22S U16558 ( .A1(n19601), .A2(n13887), .B1(n20441), .B2(n22930), .O(
        n19556) );
  AOI22S U16559 ( .A1(n19601), .A2(n21225), .B1(n20470), .B2(n22930), .O(
        n19536) );
  AOI22S U16560 ( .A1(n19601), .A2(n22932), .B1(n19634), .B2(n22930), .O(
        n19516) );
  AOI22S U16561 ( .A1(n20366), .A2(n22920), .B1(n19939), .B2(n22930), .O(
        n19476) );
  MOAI1 U16562 ( .A1(n21362), .A2(n21361), .B1(n21360), .B2(n21359), .O(n21375) );
  AN2S U16563 ( .I1(n13920), .I2(n13921), .O(n13917) );
  AN2S U16564 ( .I1(n21589), .I2(n21578), .O(n13918) );
  OR2S U16565 ( .I1(n23464), .I2(n23463), .O(n13919) );
  INV1S U16566 ( .I(n21561), .O(n21560) );
  OAI112H U16567 ( .C1(n13817), .C2(n19438), .A1(n18857), .B1(n22938), .O(
        n28527) );
  XOR2HS U16568 ( .I1(rgb_value[8]), .I2(n23462), .O(n13920) );
  XOR2HS U16569 ( .I1(n23453), .I2(n23452), .O(n13921) );
  AN2S U16570 ( .I1(n23454), .I2(n23445), .O(n13922) );
  OR2 U16571 ( .I1(n24769), .I2(n21416), .O(n13923) );
  OA112 U16572 ( .C1(n13817), .C2(n22941), .A1(n22939), .B1(n22938), .O(n13925) );
  OAI112H U16573 ( .C1(n20947), .C2(n19438), .A1(n19437), .B1(n22916), .O(
        n23839) );
  MXL2HS U16574 ( .A(n19494), .B(n20396), .S(n21654), .OB(n21660) );
  OAI112HP U16575 ( .C1(n19503), .C2(n19612), .A1(n19502), .B1(n19501), .O(
        n22412) );
  INV1S U16576 ( .I(n22930), .O(n22941) );
  NR2 U16577 ( .I1(n22918), .I2(n13822), .O(n22930) );
  NR2 U16578 ( .I1(n21551), .I2(n21561), .O(n13926) );
  OR2 U16579 ( .I1(n14173), .I2(n14146), .O(n13927) );
  OR2S U16580 ( .I1(rgb_value[9]), .I2(n21507), .O(n13928) );
  INV2 U16581 ( .I(n15448), .O(n19483) );
  OR2S U16582 ( .I1(n21521), .I2(n21522), .O(n13930) );
  INV1S U16583 ( .I(n16758), .O(n17779) );
  BUF2 U16584 ( .I(n13845), .O(n19182) );
  BUF1S U16585 ( .I(n13845), .O(n16127) );
  BUF1 U16586 ( .I(n13845), .O(n18751) );
  INV1S U16587 ( .I(n13789), .O(n17336) );
  INV1S U16588 ( .I(n13789), .O(n16635) );
  BUF1S U16589 ( .I(n28318), .O(n28221) );
  BUF1S U16590 ( .I(n28318), .O(n28468) );
  BUF1S U16591 ( .I(n28318), .O(n29076) );
  BUF1 U16592 ( .I(n27746), .O(n27065) );
  BUF1S U16593 ( .I(n28318), .O(n28412) );
  BUF1 U16594 ( .I(n26822), .O(n26101) );
  BUF1 U16595 ( .I(n29414), .O(n29435) );
  BUF1 U16596 ( .I(n26822), .O(n25595) );
  BUF1 U16597 ( .I(n27746), .O(n24415) );
  BUF1 U16598 ( .I(n27990), .O(n26970) );
  BUF1 U16599 ( .I(n29414), .O(n28106) );
  BUF1 U16600 ( .I(n26822), .O(n25810) );
  BUF1S U16601 ( .I(n28318), .O(n29129) );
  BUF1S U16602 ( .I(n28318), .O(n28643) );
  BUF1S U16603 ( .I(n28083), .O(n27987) );
  BUF1S U16604 ( .I(n28318), .O(n27685) );
  BUF1S U16605 ( .I(n28318), .O(n26490) );
  BUF1S U16606 ( .I(n28318), .O(n27722) );
  BUF1S U16607 ( .I(n28318), .O(n27957) );
  BUF1S U16608 ( .I(n28318), .O(n27110) );
  BUF1 U16609 ( .I(n24374), .O(n28182) );
  BUF1 U16610 ( .I(n24193), .O(n28162) );
  BUF1S U16611 ( .I(n24193), .O(n25468) );
  BUF1 U16612 ( .I(n24374), .O(n28614) );
  BUF1 U16613 ( .I(n24374), .O(n28135) );
  BUF1 U16614 ( .I(n24374), .O(n29194) );
  BUF1 U16615 ( .I(n13781), .O(n28938) );
  BUF1S U16616 ( .I(n24193), .O(n27443) );
  BUF1 U16617 ( .I(n24374), .O(n29096) );
  BUF1 U16618 ( .I(n13781), .O(n28037) );
  BUF1 U16619 ( .I(n24374), .O(n28075) );
  BUF1 U16620 ( .I(n23941), .O(n29242) );
  BUF1 U16621 ( .I(n24193), .O(n28433) );
  BUF1 U16622 ( .I(n23941), .O(n25859) );
  BUF1 U16623 ( .I(n13781), .O(n28343) );
  BUF1 U16624 ( .I(n24374), .O(n27735) );
  MXL2HS U16625 ( .A(n21641), .B(n20386), .S(n21654), .OB(n21657) );
  AN2 U16626 ( .I1(n17456), .I2(n17455), .O(n13932) );
  INV2 U16627 ( .I(n21811), .O(n21910) );
  INV2 U16628 ( .I(n13887), .O(n15985) );
  INV2 U16629 ( .I(n22667), .O(n22713) );
  OR2 U16630 ( .I1(n13822), .I2(n16452), .O(n13933) );
  INV2 U16631 ( .I(n22054), .O(n22171) );
  OR2 U16632 ( .I1(n21081), .I2(n21601), .O(n13935) );
  OR2 U16633 ( .I1(n28528), .I2(n20535), .O(n13938) );
  AO12 U16634 ( .B1(n22927), .B2(n21259), .A1(n19452), .O(n21236) );
  XNR2HS U16635 ( .I1(img_size[4]), .I2(n16171), .O(n13939) );
  BUF1S U16636 ( .I(n28254), .O(n24434) );
  BUF1S U16637 ( .I(n28043), .O(n29257) );
  BUF1S U16638 ( .I(n28043), .O(n26091) );
  BUF1S U16639 ( .I(n28043), .O(n24808) );
  BUF1S U16640 ( .I(n28043), .O(n26504) );
  BUF1S U16641 ( .I(n28043), .O(n24890) );
  BUF1 U16642 ( .I(n28254), .O(n24946) );
  BUF1 U16643 ( .I(n28043), .O(n27919) );
  AOI112HS U16644 ( .C1(n29996), .C2(n29999), .A1(n29995), .B1(n30021), .O(
        n13940) );
  BUF1 U16645 ( .I(n14044), .O(n19715) );
  BUF2 U16646 ( .I(n14044), .O(n18201) );
  BUF1 U16647 ( .I(n19245), .O(n19024) );
  BUF1 U16648 ( .I(n19245), .O(n20109) );
  OAI12HS U16649 ( .B1(n23827), .B2(n23826), .A1(n23825), .O(n13941) );
  BUF2 U16650 ( .I(n20039), .O(n18922) );
  BUF1S U16651 ( .I(n20039), .O(n20198) );
  BUF1S U16652 ( .I(n20039), .O(n19647) );
  BUF6 U16653 ( .I(n19642), .O(n17611) );
  BUF3 U16654 ( .I(n16016), .O(n19648) );
  BUF1 U16655 ( .I(n15568), .O(n19342) );
  BUF1S U16656 ( .I(n15568), .O(n19265) );
  INV2 U16657 ( .I(n13831), .O(n20032) );
  INV2 U16658 ( .I(n13872), .O(n19343) );
  XOR2HS U16659 ( .I1(row[3]), .I2(n23867), .O(n13942) );
  AN2S U16660 ( .I1(n21053), .I2(n22923), .O(n13943) );
  OR2 U16661 ( .I1(n23811), .I2(n14250), .O(n13946) );
  OR2 U16662 ( .I1(n14075), .I2(n14173), .O(n13947) );
  INV1S U16663 ( .I(n20956), .O(n20957) );
  ND2 U16664 ( .I1(n17697), .I2(n22058), .O(n17443) );
  AOI22S U16665 ( .A1(n13823), .A2(img[1468]), .B1(n18751), .B2(img[1340]), 
        .O(n17783) );
  OR2 U16666 ( .I1(n27889), .I2(n21637), .O(n21131) );
  AOI22S U16667 ( .A1(n13786), .A2(img[1973]), .B1(n13794), .B2(img[1845]), 
        .O(n18877) );
  AN4S U16668 ( .I1(n17771), .I2(n17770), .I3(n17769), .I4(n17768), .O(n17772)
         );
  AN4S U16669 ( .I1(n17807), .I2(n17806), .I3(n17805), .I4(n17804), .O(n17808)
         );
  AN4S U16670 ( .I1(n17621), .I2(n17620), .I3(n17619), .I4(n17618), .O(n17622)
         );
  AOI22S U16671 ( .A1(n19193), .A2(img[1789]), .B1(n17827), .B2(img[1661]), 
        .O(n19014) );
  AN4S U16672 ( .I1(n19005), .I2(n19004), .I3(n19003), .I4(n19002), .O(n19006)
         );
  AN4S U16673 ( .I1(n18915), .I2(n18914), .I3(n18913), .I4(n18912), .O(n18916)
         );
  AN4S U16674 ( .I1(n16530), .I2(n16529), .I3(n16528), .I4(n16527), .O(n16536)
         );
  AOI22S U16675 ( .A1(n19641), .A2(img[943]), .B1(n13898), .B2(img[815]), .O(
        n19306) );
  AOI22S U16676 ( .A1(n17382), .A2(img[1732]), .B1(n17862), .B2(img[1604]), 
        .O(n18721) );
  INV1S U16677 ( .I(n14045), .O(n14046) );
  MOAI1S U16678 ( .A1(n18109), .A2(n30313), .B1(n15786), .B2(img[382]), .O(
        n15482) );
  MOAI1S U16679 ( .A1(n13894), .A2(n30468), .B1(n15786), .B2(img[262]), .O(
        n15426) );
  MOAI1S U16680 ( .A1(n13850), .A2(n30821), .B1(n15809), .B2(img[1885]), .O(
        n14968) );
  MOAI1S U16681 ( .A1(n15698), .A2(n30814), .B1(n15809), .B2(img[1853]), .O(
        n15020) );
  BUF1S U16682 ( .I(n20039), .O(n18548) );
  AN4S U16683 ( .I1(n17726), .I2(n17725), .I3(n17724), .I4(n17723), .O(n17727)
         );
  AN4S U16684 ( .I1(n17844), .I2(n17843), .I3(n17842), .I4(n17841), .O(n17845)
         );
  AOI22S U16685 ( .A1(n20109), .A2(img[1417]), .B1(n13798), .B2(img[1289]), 
        .O(n16813) );
  ND2 U16686 ( .I1(n17785), .I2(n17784), .O(n20523) );
  AN4S U16687 ( .I1(n16570), .I2(n16569), .I3(n16568), .I4(n16567), .O(n16576)
         );
  AOI22S U16688 ( .A1(n19036), .A2(img[1979]), .B1(n13832), .B2(img[1851]), 
        .O(n18183) );
  MOAI1S U16689 ( .A1(n14896), .A2(n31350), .B1(n15786), .B2(img[315]), .O(
        n14898) );
  MOAI1S U16690 ( .A1(n13850), .A2(n31415), .B1(n15080), .B2(img[1971]), .O(
        n14753) );
  AN4S U16691 ( .I1(n17496), .I2(n17495), .I3(n17494), .I4(n17493), .O(n17497)
         );
  AN4S U16692 ( .I1(n17604), .I2(n17603), .I3(n17602), .I4(n17601), .O(n17610)
         );
  ND2 U16693 ( .I1(n17487), .I2(n17486), .O(n20422) );
  AN4S U16694 ( .I1(n19186), .I2(n19185), .I3(n19184), .I4(n19183), .O(n19187)
         );
  AN4S U16695 ( .I1(n19100), .I2(n19099), .I3(n19098), .I4(n19097), .O(n19101)
         );
  AN4S U16696 ( .I1(n16344), .I2(n16343), .I3(n16342), .I4(n16341), .O(n16345)
         );
  AN4S U16697 ( .I1(n16282), .I2(n16281), .I3(n16280), .I4(n16279), .O(n16283)
         );
  ND2 U16698 ( .I1(n18941), .I2(n18940), .O(n20083) );
  AN4S U16699 ( .I1(n18123), .I2(n18122), .I3(n18121), .I4(n18120), .O(n18124)
         );
  AN4S U16700 ( .I1(n18017), .I2(n18016), .I3(n18015), .I4(n18014), .O(n18018)
         );
  AN4S U16701 ( .I1(n19415), .I2(n19414), .I3(n19413), .I4(n19412), .O(n19423)
         );
  AN4S U16702 ( .I1(n19294), .I2(n19293), .I3(n19292), .I4(n19291), .O(n19301)
         );
  MOAI1S U16703 ( .A1(n15631), .A2(n31967), .B1(n13879), .B2(img[476]), .O(
        n15327) );
  MOAI1S U16704 ( .A1(n15698), .A2(n31847), .B1(n15809), .B2(img[1828]), .O(
        n15223) );
  MOAI1S U16705 ( .A1(n15668), .A2(n31827), .B1(n22928), .B2(img[1988]), .O(
        n15210) );
  MOAI1S U16706 ( .A1(n15631), .A2(n31983), .B1(n13879), .B2(img[508]), .O(
        n15158) );
  AN4S U16707 ( .I1(n18744), .I2(n18743), .I3(n18742), .I4(n18741), .O(n18745)
         );
  AOI22S U16708 ( .A1(n19667), .A2(n20963), .B1(n21062), .B2(n19663), .O(
        n19688) );
  NR2 U16709 ( .I1(n15550), .I2(n15549), .O(n15553) );
  NR2 U16710 ( .I1(n15526), .I2(n15525), .O(n15529) );
  MAOI1S U16711 ( .A1(n15660), .A2(img[254]), .B1(n30303), .B2(n15780), .O(
        n15478) );
  AN4S U16712 ( .I1(n15463), .I2(n15462), .I3(n15461), .I4(n15460), .O(n15470)
         );
  NR2 U16713 ( .I1(n15120), .I2(n15119), .O(n15122) );
  NR2 U16714 ( .I1(n15091), .I2(n15090), .O(n15094) );
  MAOI1S U16715 ( .A1(n19036), .A2(img[1909]), .B1(n30878), .B2(n15698), .O(
        n15067) );
  NR2 U16716 ( .I1(n15041), .I2(n15040), .O(n15044) );
  MAOI1S U16717 ( .A1(n19709), .A2(img[477]), .B1(n30795), .B2(n15780), .O(
        n14975) );
  NR2 U16718 ( .I1(n14942), .I2(n14941), .O(n14945) );
  MOAI1S U16719 ( .A1(n13894), .A2(n31240), .B1(n15786), .B2(img[313]), .O(
        n14162) );
  AN4S U16720 ( .I1(n15005), .I2(n15004), .I3(n15003), .I4(n15002), .O(n15012)
         );
  ND2 U16721 ( .I1(n17871), .I2(n17870), .O(n20510) );
  ND2 U16722 ( .I1(n17892), .I2(n17891), .O(n20509) );
  AN4S U16723 ( .I1(n17381), .I2(n17380), .I3(n17379), .I4(n17378), .O(n17389)
         );
  AN4S U16724 ( .I1(n16863), .I2(n16862), .I3(n16861), .I4(n16860), .O(n16869)
         );
  AN4S U16725 ( .I1(n16782), .I2(n16781), .I3(n16780), .I4(n16779), .O(n16783)
         );
  INV2 U16726 ( .I(n13872), .O(n20102) );
  ND2 U16727 ( .I1(n16576), .I2(n16575), .O(n20555) );
  AN4S U16728 ( .I1(n18290), .I2(n18289), .I3(n18288), .I4(n18287), .O(n18291)
         );
  AN4S U16729 ( .I1(n18245), .I2(n18244), .I3(n18243), .I4(n18242), .O(n18251)
         );
  AN4S U16730 ( .I1(n18169), .I2(n18168), .I3(n18167), .I4(n18166), .O(n18175)
         );
  NR2 U16731 ( .I1(n14898), .I2(n14897), .O(n14901) );
  MAOI1S U16732 ( .A1(n15568), .A2(img[891]), .B1(n31353), .B2(n15780), .O(
        n14875) );
  NR2 U16733 ( .I1(n14748), .I2(n14747), .O(n14751) );
  ND2 U16734 ( .I1(n17588), .I2(n17587), .O(n20426) );
  ND2 U16735 ( .I1(n17466), .I2(n17465), .O(n20412) );
  MOAI1S U16736 ( .A1(n15780), .A2(n27688), .B1(n15786), .B2(img[331]), .O(
        n14741) );
  MOAI1S U16737 ( .A1(n15668), .A2(n31459), .B1(n15809), .B2(img[1883]), .O(
        n14767) );
  ND2 U16738 ( .I1(n17453), .I2(n17452), .O(n19634) );
  ND2 U16739 ( .I1(n19157), .I2(n19156), .O(n19988) );
  AN4S U16740 ( .I1(n16368), .I2(n16367), .I3(n16366), .I4(n16365), .O(n16369)
         );
  ND2 U16741 ( .I1(n16346), .I2(n16345), .O(n20579) );
  ND2 U16742 ( .I1(n16677), .I2(n16676), .O(n20541) );
  AN4S U16743 ( .I1(n18647), .I2(n18646), .I3(n18645), .I4(n18644), .O(n18648)
         );
  AN4S U16744 ( .I1(n18521), .I2(n18520), .I3(n18519), .I4(n18518), .O(n18522)
         );
  ND2 U16745 ( .I1(n18094), .I2(n18093), .O(n19879) );
  ND2 U16746 ( .I1(n18019), .I2(n18018), .O(n19891) );
  ND2 U16747 ( .I1(n19409), .I2(n19408), .O(n20240) );
  AN4S U16748 ( .I1(n15230), .I2(n15229), .I3(n15228), .I4(n15227), .O(n15237)
         );
  ND2 U16749 ( .I1(n18844), .I2(n18843), .O(n20138) );
  ND2 U16750 ( .I1(n18746), .I2(n18745), .O(n20149) );
  AN4S U16751 ( .I1(n15173), .I2(n15172), .I3(n15171), .I4(n15170), .O(n15180)
         );
  AOI12HS U16752 ( .B1(n19979), .B2(n20363), .A1(n13944), .O(n19981) );
  AOI22S U16753 ( .A1(n19036), .A2(img[1984]), .B1(n13832), .B2(img[1856]), 
        .O(n18369) );
  OAI22S U16754 ( .A1(n16720), .A2(n13945), .B1(n16728), .B2(n13766), .O(
        n15152) );
  MOAI1S U16755 ( .A1(n13850), .A2(n30221), .B1(n15751), .B2(img[1839]), .O(
        n15651) );
  ND3S U16756 ( .I1(n15470), .I2(n15469), .I3(n15468), .O(n16465) );
  AN4S U16757 ( .I1(n15129), .I2(n15128), .I3(n15127), .I4(n15126), .O(n15136)
         );
  ND3S U16758 ( .I1(n14945), .I2(n14944), .I3(n14943), .O(n14952) );
  MOAI1S U16759 ( .A1(n13789), .A2(n30538), .B1(n15786), .B2(img[370]), .O(
        n14393) );
  MOAI1S U16760 ( .A1(n13850), .A2(n30739), .B1(n15080), .B2(img[1954]), .O(
        n14343) );
  MOAI1S U16761 ( .A1(n15698), .A2(n31060), .B1(n15809), .B2(img[1913]), .O(
        n14071) );
  NR2 U16762 ( .I1(n14162), .I2(n14161), .O(n14165) );
  NR2 U16763 ( .I1(n14121), .I2(n14120), .O(n14124) );
  MOAI1S U16764 ( .A1(n13789), .A2(n31192), .B1(n15786), .B2(img[329]), .O(
        n14113) );
  MOAI1S U16765 ( .A1(n15113), .A2(n31707), .B1(n15786), .B2(img[296]), .O(
        n14679) );
  MOAI1S U16766 ( .A1(n16485), .A2(n17397), .B1(n16484), .B2(n18040), .O(
        n16486) );
  MOAI1S U16767 ( .A1(n15780), .A2(n31204), .B1(n15751), .B2(img[1905]), .O(
        n14059) );
  OR2 U16768 ( .I1(i_col[1]), .I2(n23592), .O(n14173) );
  BUF1S U16769 ( .I(n18040), .O(n20968) );
  AN4S U16770 ( .I1(n16913), .I2(n16912), .I3(n16911), .I4(n16910), .O(n16914)
         );
  AN4S U16771 ( .I1(n16137), .I2(n16136), .I3(n16135), .I4(n16134), .O(n16143)
         );
  AN4S U16772 ( .I1(n17872), .I2(n17908), .I3(n17911), .I4(n17910), .O(n17873)
         );
  AN4S U16773 ( .I1(n16877), .I2(n16876), .I3(n16875), .I4(n16874), .O(n16878)
         );
  ND2 U16774 ( .I1(n18304), .I2(n18303), .O(n19663) );
  AN4S U16775 ( .I1(n14913), .I2(n14912), .I3(n14911), .I4(n14910), .O(n14921)
         );
  ND3S U16776 ( .I1(n14751), .I2(n14750), .I3(n14749), .O(n14758) );
  AN4S U16777 ( .I1(n14838), .I2(n14837), .I3(n14836), .I4(n14835), .O(n14845)
         );
  ND2 U16778 ( .I1(n16411), .I2(n16410), .O(n20581) );
  AN4S U16779 ( .I1(n18956), .I2(n18955), .I3(n18954), .I4(n18953), .O(n19049)
         );
  ND2 U16780 ( .I1(n18588), .I2(n18587), .O(n19753) );
  MOAI1S U16781 ( .A1(n17417), .A2(n17679), .B1(n17399), .B2(n20613), .O(
        n14490) );
  AN4S U16782 ( .I1(n19396), .I2(n19395), .I3(n19394), .I4(n19393), .O(n19397)
         );
  AN4S U16783 ( .I1(n15293), .I2(n15292), .I3(n15291), .I4(n15290), .O(n15300)
         );
  ND3S U16784 ( .I1(n15167), .I2(n15166), .I3(n15165), .O(n15168) );
  ND3S U16785 ( .I1(n20296), .I2(n20295), .I3(n20294), .O(n20297) );
  AN4S U16786 ( .I1(n20190), .I2(n20248), .I3(n20189), .I4(n20188), .O(n20210)
         );
  AN4S U16787 ( .I1(n18501), .I2(n18500), .I3(n18499), .I4(n18498), .O(n18502)
         );
  AN4S U16788 ( .I1(n18433), .I2(n18432), .I3(n18431), .I4(n18430), .O(n18434)
         );
  AN4S U16789 ( .I1(n18445), .I2(n18444), .I3(n18443), .I4(n18442), .O(n18446)
         );
  NR2 U16790 ( .I1(n15153), .I2(n15152), .O(n15154) );
  NR2 U16791 ( .I1(n15761), .I2(n15760), .O(n15764) );
  NR2 U16792 ( .I1(n15734), .I2(n15733), .O(n15737) );
  MOAI1S U16793 ( .A1(n15698), .A2(n30150), .B1(n15751), .B2(img[1895]), .O(
        n15729) );
  AN4S U16794 ( .I1(n15695), .I2(n15694), .I3(n15693), .I4(n15692), .O(n15703)
         );
  MOAI1S U16795 ( .A1(n15698), .A2(n30149), .B1(n15751), .B2(img[1887]), .O(
        n15617) );
  ND3S U16796 ( .I1(n15548), .I2(n15547), .I3(n15546), .O(n16481) );
  ND3S U16797 ( .I1(n15112), .I2(n15111), .I3(n15110), .O(n16727) );
  NR2 U16798 ( .I1(n14462), .I2(n14461), .O(n14465) );
  MAOI1S U16799 ( .A1(n13896), .A2(img[458]), .B1(n30549), .B2(n15780), .O(
        n14420) );
  ND3S U16800 ( .I1(n14402), .I2(n14401), .I3(n14400), .O(n14403) );
  AN4S U16801 ( .I1(n14363), .I2(n14362), .I3(n14361), .I4(n14360), .O(n14370)
         );
  MOAI1S U16802 ( .A1(n15668), .A2(n30733), .B1(n15751), .B2(img[1882]), .O(
        n14309) );
  NR2 U16803 ( .I1(n14288), .I2(n14287), .O(n14291) );
  ND3S U16804 ( .I1(n14165), .I2(n14164), .I3(n14163), .O(n14172) );
  MAOI1S U16805 ( .A1(n19023), .A2(img[1912]), .B1(n31544), .B2(n15698), .O(
        n14509) );
  NR2 U16806 ( .I1(n16487), .I2(n16486), .O(n16496) );
  MOAI1S U16807 ( .A1(n17933), .A2(n19462), .B1(n17932), .B2(n17931), .O(
        n17934) );
  AN4S U16808 ( .I1(n14219), .I2(n14218), .I3(n14217), .I4(n14216), .O(n14226)
         );
  MOAI1S U16809 ( .A1(n15765), .A2(n31534), .B1(n13797), .B2(img[736]), .O(
        n14581) );
  AN4S U16810 ( .I1(n14591), .I2(n14590), .I3(n14589), .I4(n14588), .O(n14598)
         );
  MOAI1S U16811 ( .A1(n15668), .A2(n31594), .B1(n15809), .B2(img[1872]), .O(
        n14626) );
  NR2 U16812 ( .I1(n14631), .I2(n14630), .O(n14634) );
  AN4S U16813 ( .I1(n17123), .I2(n17122), .I3(n17121), .I4(n17120), .O(n17124)
         );
  ND3S U16814 ( .I1(n23875), .I2(n23874), .I3(n28540), .O(n23876) );
  ND3S U16815 ( .I1(n26018), .I2(n28555), .I3(n26017), .O(n26019) );
  NR2 U16816 ( .I1(n14857), .I2(n14856), .O(n17675) );
  ND2 U16817 ( .I1(n18629), .I2(n18628), .O(n20324) );
  MOAI1 U16818 ( .A1(n17916), .A2(n13844), .B1(n17915), .B2(n13847), .O(n15253) );
  ND3 U16819 ( .I1(n19699), .I2(n19698), .I3(n19697), .O(n19706) );
  ND2 U16820 ( .I1(n18359), .I2(n18358), .O(n19839) );
  AOI13HS U16821 ( .B1(n15156), .B2(n15155), .B3(n15154), .A1(n20969), .O(
        n19495) );
  OR2 U16822 ( .I1(i_col[0]), .I2(i_col[1]), .O(n14251) );
  ND3S U16823 ( .I1(n15742), .I2(n15741), .I3(n15740), .O(n15743) );
  AN4S U16824 ( .I1(n15642), .I2(n15641), .I3(n15640), .I4(n15639), .O(n15649)
         );
  AN4S U16825 ( .I1(n14453), .I2(n14452), .I3(n14451), .I4(n14450), .O(n14460)
         );
  ND3S U16826 ( .I1(n14397), .I2(n14396), .I3(n14395), .O(n14398) );
  NR2 U16827 ( .I1(n14306), .I2(n14305), .O(n14313) );
  NR2 U16828 ( .I1(n14102), .I2(n14101), .O(n16935) );
  INV1S U16829 ( .I(n14251), .O(n14278) );
  ND3S U16830 ( .I1(n16496), .I2(n16495), .I3(n16494), .O(n16497) );
  NR3 U16831 ( .I1(n17927), .I2(n17926), .I3(n17925), .O(n17945) );
  MOAI1S U16832 ( .A1(n16946), .A2(n17658), .B1(n16945), .B2(n20263), .O(
        n16950) );
  AN4S U16833 ( .I1(n14580), .I2(n14579), .I3(n14578), .I4(n14577), .O(n14587)
         );
  ND3S U16834 ( .I1(n14659), .I2(n14658), .I3(n14657), .O(n14666) );
  AN4S U16835 ( .I1(n19449), .I2(n19448), .I3(n19447), .I4(n19446), .O(n19450)
         );
  AOI12HS U16836 ( .B1(n17949), .B2(n19533), .A1(n17948), .O(n17950) );
  ND2 U16837 ( .I1(n17049), .I2(n17048), .O(n21060) );
  ND2 U16838 ( .I1(n16979), .I2(n16978), .O(n21044) );
  NR2 U16839 ( .I1(n17661), .I2(n17660), .O(n17668) );
  INV1S U16840 ( .I(n26013), .O(n21597) );
  INV1S U16841 ( .I(i_col[1]), .O(n23788) );
  ND3S U16842 ( .I1(n15831), .I2(n15830), .I3(n15829), .O(n15832) );
  NR2 U16843 ( .I1(n14708), .I2(n14707), .O(n14712) );
  ND3S U16844 ( .I1(n15732), .I2(n15731), .I3(n15730), .O(n16247) );
  NR2 U16845 ( .I1(n15089), .I2(n15088), .O(n15140) );
  NR2 U16846 ( .I1(n14565), .I2(n14564), .O(n17172) );
  ND3 U16847 ( .I1(n14587), .I2(n14586), .I3(n14585), .O(n17178) );
  ND3S U16848 ( .I1(n19455), .I2(n19454), .I3(n19453), .O(n19456) );
  ND3P U16849 ( .I1(n17960), .I2(n17959), .I3(n17958), .O(n21808) );
  FA1S U16850 ( .A(rgb_value[6]), .B(rgb_value[22]), .CI(rgb_value[14]), .CO(
        n21521), .S(n21520) );
  ND3S U16851 ( .I1(n24781), .I2(n24780), .I3(n24779), .O(n24786) );
  ND3S U16852 ( .I1(n25398), .I2(n25397), .I3(n25396), .O(n25414) );
  ND3S U16853 ( .I1(n27280), .I2(n27279), .I3(n27278), .O(n27281) );
  ND3S U16854 ( .I1(n17668), .I2(n17667), .I3(n17666), .O(n17685) );
  ND2P U16855 ( .I1(n22053), .I2(n20809), .O(n21449) );
  INV1S U16856 ( .I(n23185), .O(n23294) );
  ND3S U16857 ( .I1(n15578), .I2(n15577), .I3(n15576), .O(n15579) );
  OA22 U16858 ( .A1(n20421), .A2(n17165), .B1(n17164), .B2(n17656), .O(n17169)
         );
  INV1S U16859 ( .I(n22416), .O(n22461) );
  INV1S U16860 ( .I(n21808), .O(n21914) );
  INV1S U16861 ( .I(img_size[4]), .O(n23589) );
  NR2 U16862 ( .I1(n21517), .I2(n21518), .O(n21540) );
  NR2 U16863 ( .I1(n21511), .I2(n21512), .O(n21584) );
  ND3S U16864 ( .I1(n27912), .I2(n27911), .I3(n27910), .O(n27913) );
  ND2P U16865 ( .I1(n21805), .I2(n20809), .O(n21595) );
  OAI12HS U16866 ( .B1(n29513), .B2(n13844), .A1(n15594), .O(n20605) );
  INV1S U16867 ( .I(n21660), .O(n22322) );
  OA112S U16868 ( .C1(n23763), .C2(n24030), .A1(n23762), .B1(n23761), .O(
        n23764) );
  ND3S U16869 ( .I1(n29867), .I2(n29866), .I3(n29865), .O(n29868) );
  ND2P U16870 ( .I1(n21803), .I2(n20809), .O(n21467) );
  FA1S U16871 ( .A(n15874), .B(n15873), .CI(n15872), .CO(n15881), .S(n15896)
         );
  OR2P U16872 ( .I1(n13844), .I2(n13822), .O(n18134) );
  FA1S U16873 ( .A(n22338), .B(n22337), .CI(n22336), .CO(n22356), .S(n22371)
         );
  FA1S U16874 ( .A(n22347), .B(n22346), .CI(n22345), .CO(n22362), .S(n22372)
         );
  ND3S U16875 ( .I1(n29897), .I2(n23599), .I3(n30032), .O(n29967) );
  NR2 U16876 ( .I1(n24692), .I2(n23975), .O(n24203) );
  NR2 U16877 ( .I1(n24692), .I2(n24250), .O(n24238) );
  NR2 U16878 ( .I1(n24463), .I2(n24716), .O(n24367) );
  NR2 U16879 ( .I1(n24692), .I2(n24543), .O(n24546) );
  NR2 U16880 ( .I1(n24345), .I2(n24304), .O(n24289) );
  BUF6 U16881 ( .I(n27170), .O(n27070) );
  NR2P U16882 ( .I1(n24013), .I2(n24111), .O(n24250) );
  NR2 U16883 ( .I1(i_col[3]), .I2(n23792), .O(n23835) );
  NR2 U16884 ( .I1(n21632), .I2(n21631), .O(n15915) );
  FA1S U16885 ( .A(n15861), .B(n15860), .CI(n15859), .CO(n15843), .S(n15917)
         );
  NR2 U16886 ( .I1(n23501), .I2(n23502), .O(n23503) );
  FA1S U16887 ( .A(n15964), .B(n15963), .CI(n15962), .CO(n15994), .S(n15976)
         );
  FA1S U16888 ( .A(n22366), .B(n22365), .CI(n22364), .CO(n22361), .S(n22396)
         );
  ND3S U16889 ( .I1(n23774), .I2(n23773), .I3(n23772), .O(n23783) );
  INV1S U16890 ( .I(n21571), .O(n21563) );
  FA1S U16891 ( .A(n15842), .B(n15841), .CI(n15840), .CO(n21774), .S(n21781)
         );
  MOAI1 U16892 ( .A1(n23504), .A2(n23503), .B1(n23502), .B2(n23501), .O(n23519) );
  ND3S U16893 ( .I1(n23730), .I2(n23729), .I3(n23774), .O(n23739) );
  TIE1 U16894 ( .O(n11230) );
  XOR2HS U16895 ( .I1(n23900), .I2(img_size[3]), .O(n23859) );
  OR2 U16896 ( .I1(img_size[0]), .I2(img_size[1]), .O(n23973) );
  INV1S U16897 ( .I(n23973), .O(n24332) );
  NR2 U16898 ( .I1(img_size[3]), .I2(n23589), .O(n13948) );
  INV1S U16899 ( .I(img_size[5]), .O(n23665) );
  OAI12HS U16900 ( .B1(n13949), .B2(n24698), .A1(n23897), .O(n24031) );
  INV1S U16901 ( .I(addr[1]), .O(n30004) );
  INV1S U16902 ( .I(n23897), .O(n24701) );
  MOAI1S U16903 ( .A1(addr[0]), .A2(addr[2]), .B1(addr[0]), .B2(addr[3]), .O(
        n13952) );
  NR2 U16904 ( .I1(addr[7]), .I2(addr[6]), .O(n23618) );
  NR2 U16905 ( .I1(n23618), .I2(n24701), .O(n13951) );
  AN4B1S U16906 ( .I1(n13954), .I2(n13953), .I3(n13952), .B1(n13951), .O(
        n13956) );
  MOAI1S U16907 ( .A1(addr[3]), .A2(addr[1]), .B1(n24031), .B2(addr[2]), .O(
        n13955) );
  INV1S U16908 ( .I(n24698), .O(n23898) );
  NR2 U16909 ( .I1(addr[5]), .I2(addr[4]), .O(n23619) );
  MOAI1S U16910 ( .A1(n23923), .A2(n23619), .B1(n23923), .B2(n23560), .O(
        n13957) );
  NR2 U16911 ( .I1(n13958), .I2(n13957), .O(n30026) );
  INV2 U16912 ( .I(act_ptr[2]), .O(n23642) );
  ND2S U16913 ( .I1(n13986), .I2(act[1]), .O(n13961) );
  ND2S U16914 ( .I1(n13987), .I2(act[13]), .O(n13960) );
  ND3S U16915 ( .I1(n13961), .I2(n13960), .I3(act_ptr[0]), .O(n13968) );
  INV1S U16916 ( .I(n13989), .O(n23641) );
  INV1S U16917 ( .I(act[7]), .O(n13962) );
  MOAI1 U16918 ( .A1(n23641), .A2(n13962), .B1(n13988), .B2(act[19]), .O(
        n13967) );
  AOI22S U16919 ( .A1(n13987), .A2(act[16]), .B1(n13986), .B2(act[4]), .O(
        n13965) );
  AOI12HS U16920 ( .B1(n13988), .B2(act[22]), .A1(act_ptr[0]), .O(n13964) );
  INV1S U16921 ( .I(n23852), .O(n13996) );
  INV1S U16922 ( .I(act[15]), .O(n13969) );
  INV2 U16923 ( .I(n13987), .O(n23639) );
  INV1S U16924 ( .I(n13988), .O(n13984) );
  INV1S U16925 ( .I(act[21]), .O(n23884) );
  OAI22S U16926 ( .A1(n13969), .A2(n23639), .B1(n13984), .B2(n23884), .O(
        n13973) );
  ND2S U16927 ( .I1(n13989), .I2(act[9]), .O(n13970) );
  NR2 U16928 ( .I1(n13973), .I2(n13972), .O(n13980) );
  INV1S U16929 ( .I(act[12]), .O(n13974) );
  MOAI1 U16930 ( .A1(n23639), .A2(n13974), .B1(n13988), .B2(act[18]), .O(
        n13978) );
  ND2S U16931 ( .I1(n13986), .I2(act[0]), .O(n13976) );
  ND2S U16932 ( .I1(n13989), .I2(act[6]), .O(n13975) );
  NR2 U16933 ( .I1(n13978), .I2(n13977), .O(n13979) );
  NR2P U16934 ( .I1(n13980), .I2(n13979), .O(n23895) );
  ND2S U16935 ( .I1(n13989), .I2(act[8]), .O(n13981) );
  INV1S U16936 ( .I(act[14]), .O(n13985) );
  INV1S U16937 ( .I(act[20]), .O(n13983) );
  OAI22S U16938 ( .A1(n13985), .A2(n23639), .B1(n13984), .B2(n13983), .O(
        n13994) );
  AOI22S U16939 ( .A1(n13987), .A2(act[17]), .B1(n13986), .B2(act[5]), .O(
        n13992) );
  AOI12HS U16940 ( .B1(n13988), .B2(act[23]), .A1(act_ptr[0]), .O(n13991) );
  OR2P U16941 ( .I1(n23851), .I2(n23852), .O(n14017) );
  OAI222S U16942 ( .A1(n23919), .A2(n23607), .B1(n13822), .B2(n24701), .C1(
        n14017), .C2(n23923), .O(n13997) );
  XNR2HS U16943 ( .I1(cal_cnt[4]), .I2(n13997), .O(n14010) );
  OAI22S U16944 ( .A1(n14017), .A2(n23919), .B1(n23607), .B2(n23897), .O(
        n13998) );
  XNR2HS U16945 ( .I1(cal_cnt[6]), .I2(n13998), .O(n14009) );
  NR2 U16946 ( .I1(n23897), .I2(n14017), .O(n14001) );
  OAI12HS U16947 ( .B1(n23895), .B2(cal_cnt[5]), .A1(n14001), .O(n14000) );
  INV12 U16948 ( .I(n13822), .O(n20809) );
  AOI22S U16949 ( .A1(cal_cnt[8]), .A2(n14000), .B1(n13999), .B2(cal_cnt[5]), 
        .O(n14008) );
  NR2 U16950 ( .I1(cal_cnt[0]), .I2(cal_cnt[1]), .O(n29971) );
  INV1S U16951 ( .I(n14001), .O(n14002) );
  NR2 U16952 ( .I1(cal_cnt[8]), .I2(n14002), .O(n14003) );
  NR3 U16953 ( .I1(cal_cnt[7]), .I2(cal_cnt[2]), .I3(n14003), .O(n14006) );
  NR2 U16954 ( .I1(n23923), .I2(n13822), .O(n14004) );
  XNR2HS U16955 ( .I1(cal_cnt[3]), .I2(n14004), .O(n14005) );
  AN4B1S U16956 ( .I1(n14010), .I2(n14009), .I3(n14008), .B1(n14007), .O(
        n14021) );
  NR2 U16957 ( .I1(n14012), .I2(n23565), .O(n23691) );
  NR2 U16958 ( .I1(n14029), .I2(c_s[1]), .O(n21501) );
  INV1S U16959 ( .I(n21501), .O(n23694) );
  INV1S U16960 ( .I(n29910), .O(n31997) );
  NR2 U16961 ( .I1(n23694), .I2(n14013), .O(n14028) );
  INV1S U16962 ( .I(n23691), .O(n14014) );
  INV1S U16963 ( .I(n23561), .O(n14026) );
  ND2S U16964 ( .I1(act[18]), .I2(act[19]), .O(n14015) );
  NR2 U16965 ( .I1(n14015), .I2(c_s[0]), .O(n14016) );
  ND3S U16966 ( .I1(n14016), .I2(act[20]), .I3(act_delay2), .O(n14020) );
  INV1S U16967 ( .I(n14017), .O(n14018) );
  NR2 U16968 ( .I1(c_s[0]), .I2(n23565), .O(n29969) );
  ND3S U16969 ( .I1(n14018), .I2(n23895), .I3(n29969), .O(n14019) );
  OAI112HS U16970 ( .C1(n23694), .C2(n14020), .A1(n14019), .B1(n23682), .O(
        n14025) );
  INV1S U16971 ( .I(set_cnt[0]), .O(n29996) );
  ND3S U16972 ( .I1(n14021), .I2(set_cnt[3]), .I3(n29996), .O(n14023) );
  NR3 U16973 ( .I1(n14026), .I2(n14025), .I3(n14024), .O(n14027) );
  OAI12HS U16974 ( .B1(in_valid), .B2(N25894), .A1(n14027), .O(n23586) );
  INV1S U16975 ( .I(n29969), .O(n29991) );
  ND2P U16976 ( .I1(in_valid), .I2(n14029), .O(n23571) );
  INV1S U16977 ( .I(c_s[0]), .O(n14030) );
  NR2 U16978 ( .I1(act_delay2), .I2(n23572), .O(n14031) );
  OA222 U16979 ( .A1(n29962), .A2(n29991), .B1(n23571), .B2(c_s[1]), .C1(
        n14032), .C2(n14031), .O(n23587) );
  INV1S U16980 ( .I(template_store[45]), .O(n21728) );
  ND2F U16981 ( .I1(i_row[1]), .I2(i_row[0]), .O(n23623) );
  NR2F U16982 ( .I1(n14033), .I2(n23623), .O(n17886) );
  OR2T U16983 ( .I1(i_row[2]), .I2(n23823), .O(n14047) );
  AOI22S U16984 ( .A1(n17793), .A2(img[113]), .B1(n15506), .B2(img[625]), .O(
        n14042) );
  OR2T U16985 ( .I1(i_row[0]), .I2(i_row[1]), .O(n23624) );
  OR2T U16986 ( .I1(i_row[1]), .I2(n23824), .O(n14058) );
  INV4 U16987 ( .I(n15786), .O(n15631) );
  INV8 U16988 ( .I(n15631), .O(n15537) );
  AOI22S U16989 ( .A1(n13895), .A2(img[497]), .B1(n15537), .B2(img[369]), .O(
        n14041) );
  ND2P U16990 ( .I1(n23824), .I2(i_row[3]), .O(n14035) );
  NR2F U16991 ( .I1(n14035), .I2(n23827), .O(n19642) );
  INV2 U16992 ( .I(n19642), .O(n14036) );
  INV6 U16993 ( .I(n14036), .O(n15660) );
  NR2T U16994 ( .I1(i_row[3]), .I2(n14037), .O(n14054) );
  INV1S U16995 ( .I(n14054), .O(n14038) );
  NR2T U16996 ( .I1(n14058), .I2(n14038), .O(n16364) );
  AOI22S U16997 ( .A1(n15660), .A2(img[241]), .B1(n13854), .B2(img[1393]), .O(
        n14040) );
  OR2T U16998 ( .I1(i_row[3]), .I2(i_row[0]), .O(n14052) );
  NR2F U16999 ( .I1(n14052), .I2(n23827), .O(n17885) );
  AOI22S U17000 ( .A1(n15800), .A2(img[1265]), .B1(n13885), .B2(img[881]), .O(
        n14039) );
  AN4S U17001 ( .I1(n14042), .I2(n14041), .I3(n14040), .I4(n14039), .O(n14063)
         );
  NR2P U17002 ( .I1(i_row[3]), .I2(i_row[2]), .O(n14056) );
  INV4CK U17003 ( .I(n13842), .O(n15698) );
  NR2T U17004 ( .I1(n23624), .I2(n14047), .O(n14111) );
  MOAI1S U17005 ( .A1(n15698), .A2(n31165), .B1(n15653), .B2(img[1009]), .O(
        n14049) );
  MOAI1S U17006 ( .A1(n15765), .A2(n31157), .B1(n13797), .B2(img[753]), .O(
        n14048) );
  NR2 U17007 ( .I1(n14049), .I2(n14048), .O(n14062) );
  OR2P U17008 ( .I1(i_row[2]), .I2(i_row[1]), .O(n14051) );
  NR2F U17009 ( .I1(n14052), .I2(n14051), .O(n22928) );
  INV6 U17010 ( .I(n14053), .O(n15080) );
  MOAI1S U17011 ( .A1(n13850), .A2(n31210), .B1(n15080), .B2(img[2033]), .O(
        n14060) );
  INV2 U17012 ( .I(n23624), .O(n14055) );
  OR2T U17013 ( .I1(n14058), .I2(n14057), .O(n14077) );
  NR2 U17014 ( .I1(n14060), .I2(n14059), .O(n14061) );
  ND3 U17015 ( .I1(n14063), .I2(n14062), .I3(n14061), .O(n16938) );
  INV1S U17016 ( .I(n16938), .O(n14076) );
  INV2 U17017 ( .I(i_col[3]), .O(n23794) );
  ND3S U17018 ( .I1(n23794), .I2(n23792), .I3(i_col[1]), .O(n14227) );
  AOI22S U17019 ( .A1(n13860), .A2(img[1017]), .B1(n15660), .B2(img[249]), .O(
        n14067) );
  AOI22S U17020 ( .A1(n15799), .A2(img[505]), .B1(n15537), .B2(img[377]), .O(
        n14066) );
  AOI22S U17021 ( .A1(n15800), .A2(img[1273]), .B1(n18298), .B2(img[1401]), 
        .O(n14065) );
  AOI22S U17022 ( .A1(n13801), .A2(img[121]), .B1(n15506), .B2(img[633]), .O(
        n14064) );
  AN4S U17023 ( .I1(n14067), .I2(n14066), .I3(n14065), .I4(n14064), .O(n14074)
         );
  MOAI1S U17024 ( .A1(n13850), .A2(n31064), .B1(n15080), .B2(img[2041]), .O(
        n14069) );
  MOAI1S U17025 ( .A1(n15765), .A2(n31052), .B1(n13898), .B2(img[761]), .O(
        n14068) );
  NR2 U17026 ( .I1(n14069), .I2(n14068), .O(n14073) );
  MOAI1S U17027 ( .A1(n15780), .A2(n31032), .B1(n13884), .B2(img[889]), .O(
        n14070) );
  NR2 U17028 ( .I1(n14071), .I2(n14070), .O(n14072) );
  ND3 U17029 ( .I1(n14074), .I2(n14073), .I3(n14072), .O(n16947) );
  INV1 U17030 ( .I(i_col[0]), .O(n23592) );
  MOAI1S U17031 ( .A1(n13850), .A2(n31207), .B1(n15080), .B2(img[1969]), .O(
        n14079) );
  MOAI1S U17032 ( .A1(n18109), .A2(n31146), .B1(n13884), .B2(img[817]), .O(
        n14078) );
  NR2 U17033 ( .I1(n14079), .I2(n14078), .O(n14082) );
  AOI22S U17034 ( .A1(n13898), .A2(img[689]), .B1(n15652), .B2(img[1713]), .O(
        n14081) );
  AOI22S U17035 ( .A1(n13858), .A2(img[433]), .B1(n15537), .B2(img[305]), .O(
        n14080) );
  ND3S U17036 ( .I1(n14082), .I2(n14081), .I3(n14080), .O(n14089) );
  INV2 U17037 ( .I(n13840), .O(n15657) );
  MOAI1S U17038 ( .A1(n15674), .A2(n31215), .B1(n15657), .B2(img[561]), .O(
        n14084) );
  INV2 U17039 ( .I(n13931), .O(n15668) );
  OAI22S U17040 ( .A1(n15698), .A2(n31162), .B1(n15668), .B2(n31201), .O(
        n14083) );
  NR2 U17041 ( .I1(n14084), .I2(n14083), .O(n14087) );
  AOI22S U17042 ( .A1(n13880), .A2(img[945]), .B1(n15660), .B2(img[177]), .O(
        n14086) );
  AOI22S U17043 ( .A1(n15800), .A2(img[1201]), .B1(n13854), .B2(img[1329]), 
        .O(n14085) );
  ND3S U17044 ( .I1(n14087), .I2(n14086), .I3(n14085), .O(n14088) );
  OR2P U17045 ( .I1(i_col[2]), .I2(n23794), .O(n14200) );
  INV2 U17046 ( .I(n14200), .O(n23834) );
  NR2 U17047 ( .I1(i_col[0]), .I2(n23788), .O(n14145) );
  MOAI1S U17048 ( .A1(n13850), .A2(n31209), .B1(n15080), .B2(img[1929]), .O(
        n14091) );
  MOAI1S U17049 ( .A1(n15765), .A2(n31156), .B1(n13837), .B2(img[649]), .O(
        n14090) );
  NR2 U17050 ( .I1(n14091), .I2(n14090), .O(n14095) );
  AOI22S U17051 ( .A1(n13858), .A2(img[393]), .B1(n13845), .B2(img[1417]), .O(
        n14094) );
  INV4CK U17052 ( .I(n14092), .O(n15773) );
  AOI22S U17053 ( .A1(n13892), .A2(img[905]), .B1(n15773), .B2(img[137]), .O(
        n14093) );
  ND3S U17054 ( .I1(n14095), .I2(n14094), .I3(n14093), .O(n14102) );
  MOAI1S U17055 ( .A1(n15698), .A2(n31164), .B1(n15786), .B2(img[265]), .O(
        n14097) );
  MOAI1S U17056 ( .A1(n18109), .A2(n31148), .B1(n15568), .B2(img[777]), .O(
        n14096) );
  NR2 U17057 ( .I1(n14097), .I2(n14096), .O(n14100) );
  AOI22S U17058 ( .A1(n13802), .A2(img[1161]), .B1(n13853), .B2(img[1289]), 
        .O(n14099) );
  AOI22S U17059 ( .A1(n14909), .A2(img[9]), .B1(n15506), .B2(img[521]), .O(
        n14098) );
  ND3 U17060 ( .I1(n14100), .I2(n14099), .I3(n14098), .O(n14101) );
  ND2S U17061 ( .I1(i_col[1]), .I2(i_col[0]), .O(n23811) );
  ND2 U17062 ( .I1(i_col[3]), .I2(i_col[2]), .O(n14250) );
  OAI22S U17063 ( .A1(n16946), .A2(n16468), .B1(n16935), .B2(n13946), .O(
        n14103) );
  NR2 U17064 ( .I1(n14104), .I2(n14103), .O(n14160) );
  INV1S U17065 ( .I(n23811), .O(n14105) );
  BUF1 U17066 ( .I(n18040), .O(n20629) );
  MOAI1S U17067 ( .A1(n15765), .A2(n31155), .B1(n13898), .B2(img[713]), .O(
        n14109) );
  AOI22S U17068 ( .A1(n13895), .A2(img[457]), .B1(n15568), .B2(img[841]), .O(
        n14107) );
  ND2S U17069 ( .I1(n15773), .I2(img[201]), .O(n14106) );
  OAI112HS U17070 ( .C1(n15668), .C2(n31202), .A1(n14107), .B1(n14106), .O(
        n14108) );
  NR3 U17071 ( .I1(n14110), .I2(n14109), .I3(n14108), .O(n14119) );
  MOAI1S U17072 ( .A1(n19648), .A2(n31218), .B1(n14909), .B2(img[73]), .O(
        n14114) );
  NR2 U17073 ( .I1(n14114), .I2(n14113), .O(n14118) );
  MOAI1S U17074 ( .A1(n15698), .A2(n31163), .B1(n15751), .B2(img[1865]), .O(
        n14116) );
  MOAI1S U17075 ( .A1(n13838), .A2(n31183), .B1(n15657), .B2(img[585]), .O(
        n14115) );
  NR2 U17076 ( .I1(n14116), .I2(n14115), .O(n14117) );
  ND3 U17077 ( .I1(n14119), .I2(n14118), .I3(n14117), .O(n16932) );
  MOAI1S U17078 ( .A1(n19648), .A2(n31109), .B1(n19642), .B2(img[153]), .O(
        n14120) );
  AOI22S U17079 ( .A1(n18909), .A2(img[1177]), .B1(n13853), .B2(img[1305]), 
        .O(n14123) );
  AOI22S U17080 ( .A1(n17864), .A2(img[25]), .B1(n15506), .B2(img[537]), .O(
        n14122) );
  AOI22S U17081 ( .A1(n13865), .A2(img[1817]), .B1(n15630), .B2(img[1561]), 
        .O(n14129) );
  MOAI1S U17082 ( .A1(n13850), .A2(n31100), .B1(n15080), .B2(img[1945]), .O(
        n14126) );
  MOAI1S U17083 ( .A1(n15765), .A2(n31048), .B1(n13837), .B2(img[665]), .O(
        n14125) );
  NR2 U17084 ( .I1(n14126), .I2(n14125), .O(n14128) );
  AOI22S U17085 ( .A1(n13884), .A2(img[793]), .B1(n13845), .B2(img[1433]), .O(
        n14127) );
  ND3S U17086 ( .I1(n14129), .I2(n14128), .I3(n14127), .O(n14130) );
  NR2 U17087 ( .I1(n14131), .I2(n14130), .O(n14262) );
  INV1S U17088 ( .I(n14262), .O(n16941) );
  INV1S U17089 ( .I(n14250), .O(n14133) );
  INV1S U17090 ( .I(n14173), .O(n14132) );
  AOI22S U17091 ( .A1(n20629), .A2(n16932), .B1(n16941), .B2(n17762), .O(
        n14159) );
  AOI22S U17092 ( .A1(n15653), .A2(img[977]), .B1(n15773), .B2(img[209]), .O(
        n14137) );
  AOI22S U17093 ( .A1(n18262), .A2(img[465]), .B1(n19710), .B2(img[337]), .O(
        n14136) );
  AOI22S U17094 ( .A1(n15800), .A2(img[1233]), .B1(n13853), .B2(img[1361]), 
        .O(n14135) );
  AOI22S U17095 ( .A1(n13801), .A2(img[81]), .B1(n15506), .B2(img[593]), .O(
        n14134) );
  AN4S U17096 ( .I1(n14137), .I2(n14136), .I3(n14135), .I4(n14134), .O(n14144)
         );
  MOAI1S U17097 ( .A1(n13850), .A2(n31173), .B1(n15080), .B2(img[2001]), .O(
        n14139) );
  MOAI1S U17098 ( .A1(n15765), .A2(n31161), .B1(n13837), .B2(img[721]), .O(
        n14138) );
  NR2 U17099 ( .I1(n14139), .I2(n14138), .O(n14143) );
  MOAI1S U17100 ( .A1(n15698), .A2(n31169), .B1(n15751), .B2(img[1873]), .O(
        n14141) );
  MOAI1S U17101 ( .A1(n15668), .A2(n31142), .B1(n15568), .B2(img[849]), .O(
        n14140) );
  NR2 U17102 ( .I1(n14141), .I2(n14140), .O(n14142) );
  ND3 U17103 ( .I1(n14144), .I2(n14143), .I3(n14142), .O(n16934) );
  INV1S U17104 ( .I(n23835), .O(n14146) );
  INV1S U17105 ( .I(n14145), .O(n14213) );
  INV2 U17106 ( .I(n13929), .O(n20439) );
  AOI22S U17107 ( .A1(n19258), .A2(img[985]), .B1(n15773), .B2(img[217]), .O(
        n14150) );
  AOI22S U17108 ( .A1(n13896), .A2(img[473]), .B1(n15537), .B2(img[345]), .O(
        n14149) );
  AOI22S U17109 ( .A1(n15800), .A2(img[1241]), .B1(n13854), .B2(img[1369]), 
        .O(n14148) );
  AOI22S U17110 ( .A1(n13803), .A2(img[89]), .B1(n13785), .B2(img[601]), .O(
        n14147) );
  AN4S U17111 ( .I1(n14150), .I2(n14149), .I3(n14148), .I4(n14147), .O(n14157)
         );
  MOAI1S U17112 ( .A1(n13850), .A2(n31102), .B1(n15080), .B2(img[2009]), .O(
        n14152) );
  MOAI1S U17113 ( .A1(n15765), .A2(n31047), .B1(n13797), .B2(img[729]), .O(
        n14151) );
  NR2 U17114 ( .I1(n14152), .I2(n14151), .O(n14156) );
  MOAI1S U17115 ( .A1(n15698), .A2(n31055), .B1(n15751), .B2(img[1881]), .O(
        n14154) );
  MOAI1S U17116 ( .A1(n15668), .A2(n31095), .B1(n13884), .B2(img[857]), .O(
        n14153) );
  NR2 U17117 ( .I1(n14154), .I2(n14153), .O(n14155) );
  ND3 U17118 ( .I1(n14157), .I2(n14156), .I3(n14155), .O(n16940) );
  AOI22S U17119 ( .A1(n16934), .A2(n20439), .B1(n13791), .B2(n16940), .O(
        n14158) );
  ND3 U17120 ( .I1(n14160), .I2(n14159), .I3(n14158), .O(n14256) );
  MOAI1S U17121 ( .A1(n19648), .A2(n31234), .B1(n19642), .B2(img[185]), .O(
        n14161) );
  AOI22S U17122 ( .A1(n18548), .A2(img[1209]), .B1(n13783), .B2(img[1337]), 
        .O(n14164) );
  AOI22S U17123 ( .A1(n17864), .A2(img[57]), .B1(n15506), .B2(img[569]), .O(
        n14163) );
  AOI22S U17124 ( .A1(n13865), .A2(img[1849]), .B1(n15630), .B2(img[1593]), 
        .O(n14170) );
  MOAI1S U17125 ( .A1(n13850), .A2(n31062), .B1(n15080), .B2(img[1977]), .O(
        n14167) );
  MOAI1S U17126 ( .A1(n15765), .A2(n31050), .B1(n13797), .B2(img[697]), .O(
        n14166) );
  NR2 U17127 ( .I1(n14167), .I2(n14166), .O(n14169) );
  AOI22S U17128 ( .A1(n13784), .A2(img[825]), .B1(n13845), .B2(img[1465]), .O(
        n14168) );
  ND3S U17129 ( .I1(n14170), .I2(n14169), .I3(n14168), .O(n14171) );
  NR2 U17130 ( .I1(n14173), .I2(n14200), .O(n14174) );
  MOAI1S U17131 ( .A1(n15698), .A2(n31057), .B1(n13895), .B2(img[481]), .O(
        n14176) );
  MOAI1S U17132 ( .A1(n18141), .A2(n31069), .B1(n15657), .B2(img[609]), .O(
        n14175) );
  NR2 U17133 ( .I1(n14176), .I2(n14175), .O(n14179) );
  AOI22S U17134 ( .A1(n13893), .A2(img[993]), .B1(n13824), .B2(img[1377]), .O(
        n14178) );
  AOI22S U17135 ( .A1(n18958), .A2(img[97]), .B1(n15800), .B2(img[1249]), .O(
        n14177) );
  ND3S U17136 ( .I1(n14179), .I2(n14178), .I3(n14177), .O(n14186) );
  MOAI1S U17137 ( .A1(n13850), .A2(n31101), .B1(n15751), .B2(img[1889]), .O(
        n14181) );
  MOAI1S U17138 ( .A1(n15765), .A2(n31049), .B1(n13837), .B2(img[737]), .O(
        n14180) );
  NR2 U17139 ( .I1(n14181), .I2(n14180), .O(n14184) );
  MAOI1S U17140 ( .A1(n13885), .A2(img[865]), .B1(n31094), .B2(n15668), .O(
        n14183) );
  AOI22S U17141 ( .A1(n15537), .A2(img[353]), .B1(n15773), .B2(img[225]), .O(
        n14182) );
  ND3S U17142 ( .I1(n14184), .I2(n14183), .I3(n14182), .O(n14185) );
  ND2 U17143 ( .I1(n23835), .I2(n14278), .O(n20587) );
  OAI22S U17144 ( .A1(n16954), .A2(n15142), .B1(n16933), .B2(n20587), .O(
        n14215) );
  MOAI1S U17145 ( .A1(n13894), .A2(n31137), .B1(n13885), .B2(img[809]), .O(
        n14187) );
  NR2 U17146 ( .I1(n14188), .I2(n14187), .O(n14192) );
  AOI22S U17147 ( .A1(n13883), .A2(img[553]), .B1(n16515), .B2(img[1065]), .O(
        n14191) );
  AOI22S U17148 ( .A1(n13837), .A2(img[681]), .B1(n15652), .B2(img[1705]), .O(
        n14190) );
  ND3S U17149 ( .I1(n14192), .I2(n14191), .I3(n14190), .O(n14199) );
  MOAI1S U17150 ( .A1(n15674), .A2(n31121), .B1(n15800), .B2(img[1193]), .O(
        n14194) );
  OAI22S U17151 ( .A1(n15698), .A2(n31168), .B1(n15668), .B2(n31141), .O(
        n14193) );
  NR2 U17152 ( .I1(n14194), .I2(n14193), .O(n14197) );
  AOI22S U17153 ( .A1(n15537), .A2(img[297]), .B1(n15660), .B2(img[169]), .O(
        n14196) );
  AOI22S U17154 ( .A1(n13889), .A2(img[937]), .B1(n14392), .B2(img[1321]), .O(
        n14195) );
  ND3S U17155 ( .I1(n14197), .I2(n14196), .I3(n14195), .O(n14198) );
  NR2P U17156 ( .I1(n14199), .I2(n14198), .O(n16948) );
  NR2 U17157 ( .I1(n23811), .I2(n14200), .O(n19931) );
  INV2 U17158 ( .I(n19931), .O(n17397) );
  MOAI1S U17159 ( .A1(n19648), .A2(n31248), .B1(n19642), .B2(img[145]), .O(
        n14201) );
  NR2 U17160 ( .I1(n14202), .I2(n14201), .O(n14205) );
  AOI22S U17161 ( .A1(n13792), .A2(img[1169]), .B1(n15315), .B2(img[1297]), 
        .O(n14204) );
  AOI22S U17162 ( .A1(n13841), .A2(img[17]), .B1(n15506), .B2(img[529]), .O(
        n14203) );
  ND3S U17163 ( .I1(n14205), .I2(n14204), .I3(n14203), .O(n14212) );
  AOI22S U17164 ( .A1(n13865), .A2(img[1809]), .B1(n20109), .B2(img[1553]), 
        .O(n14210) );
  MOAI1S U17165 ( .A1(n13850), .A2(n31170), .B1(n15080), .B2(img[1937]), .O(
        n14207) );
  MOAI1S U17166 ( .A1(n15765), .A2(n31158), .B1(n13837), .B2(img[657]), .O(
        n14206) );
  NR2 U17167 ( .I1(n14207), .I2(n14206), .O(n14209) );
  AOI22S U17168 ( .A1(n19641), .A2(img[785]), .B1(n13845), .B2(img[1425]), .O(
        n14208) );
  ND3S U17169 ( .I1(n14210), .I2(n14209), .I3(n14208), .O(n14211) );
  NR2P U17170 ( .I1(n14212), .I2(n14211), .O(n16951) );
  OAI22S U17171 ( .A1(n16948), .A2(n17397), .B1(n16951), .B2(n17679), .O(
        n14214) );
  NR2 U17172 ( .I1(n14215), .I2(n14214), .O(n14254) );
  AOI22S U17173 ( .A1(n19403), .A2(img[1001]), .B1(n15660), .B2(img[233]), .O(
        n14219) );
  AOI22S U17174 ( .A1(n19709), .A2(img[489]), .B1(n15537), .B2(img[361]), .O(
        n14218) );
  AOI22S U17175 ( .A1(n15800), .A2(img[1257]), .B1(n13854), .B2(img[1385]), 
        .O(n14217) );
  AOI22S U17176 ( .A1(n13801), .A2(img[105]), .B1(n15506), .B2(img[617]), .O(
        n14216) );
  MOAI1S U17177 ( .A1(n13850), .A2(n31171), .B1(n15080), .B2(img[2025]), .O(
        n14221) );
  MOAI1S U17178 ( .A1(n15765), .A2(n31159), .B1(n13797), .B2(img[745]), .O(
        n14220) );
  NR2 U17179 ( .I1(n14221), .I2(n14220), .O(n14225) );
  MOAI1S U17180 ( .A1(n15698), .A2(n31167), .B1(n15751), .B2(img[1897]), .O(
        n14223) );
  MOAI1S U17181 ( .A1(n15780), .A2(n31140), .B1(n13885), .B2(img[873]), .O(
        n14222) );
  NR2 U17182 ( .I1(n14223), .I2(n14222), .O(n14224) );
  ND3 U17183 ( .I1(n14226), .I2(n14225), .I3(n14224), .O(n16956) );
  NR2 U17184 ( .I1(n23592), .I2(n14227), .O(n14869) );
  INV2 U17185 ( .I(n14869), .O(n14259) );
  NR2 U17186 ( .I1(i_col[2]), .I2(n14251), .O(n14257) );
  INV1S U17187 ( .I(n14257), .O(n18196) );
  AOI22S U17188 ( .A1(n15653), .A2(img[961]), .B1(n15660), .B2(img[193]), .O(
        n14231) );
  AOI22S U17189 ( .A1(n13896), .A2(img[449]), .B1(n15537), .B2(img[321]), .O(
        n14230) );
  AOI22S U17190 ( .A1(n15800), .A2(img[1217]), .B1(n15315), .B2(img[1345]), 
        .O(n14229) );
  AOI22S U17191 ( .A1(n20104), .A2(img[65]), .B1(n15506), .B2(img[577]), .O(
        n14228) );
  AN4S U17192 ( .I1(n14231), .I2(n14230), .I3(n14229), .I4(n14228), .O(n14238)
         );
  MOAI1S U17193 ( .A1(n13850), .A2(n31063), .B1(n15080), .B2(img[1985]), .O(
        n14233) );
  MOAI1S U17194 ( .A1(n15765), .A2(n31051), .B1(n13797), .B2(img[705]), .O(
        n14232) );
  NR2 U17195 ( .I1(n14233), .I2(n14232), .O(n14237) );
  MOAI1S U17196 ( .A1(n15698), .A2(n31059), .B1(n15751), .B2(img[1857]), .O(
        n14235) );
  MOAI1S U17197 ( .A1(n15780), .A2(n31031), .B1(n13885), .B2(img[833]), .O(
        n14234) );
  NR2 U17198 ( .I1(n14235), .I2(n14234), .O(n14236) );
  ND3 U17199 ( .I1(n14238), .I2(n14237), .I3(n14236), .O(n16945) );
  AOI22S U17200 ( .A1(n16956), .A2(n21062), .B1(n13843), .B2(n16945), .O(
        n14253) );
  AOI22S U17201 ( .A1(n15653), .A2(img[929]), .B1(n15773), .B2(img[161]), .O(
        n14242) );
  AOI22S U17202 ( .A1(n13895), .A2(img[417]), .B1(n13800), .B2(img[289]), .O(
        n14241) );
  AOI22S U17203 ( .A1(n15800), .A2(img[1185]), .B1(n15315), .B2(img[1313]), 
        .O(n14240) );
  AOI22S U17204 ( .A1(n17864), .A2(img[33]), .B1(n15506), .B2(img[545]), .O(
        n14239) );
  AN4S U17205 ( .I1(n14242), .I2(n14241), .I3(n14240), .I4(n14239), .O(n14249)
         );
  MOAI1S U17206 ( .A1(n13850), .A2(n31103), .B1(n15080), .B2(img[1953]), .O(
        n14244) );
  MOAI1S U17207 ( .A1(n15765), .A2(n31046), .B1(n13898), .B2(img[673]), .O(
        n14243) );
  NR2 U17208 ( .I1(n14244), .I2(n14243), .O(n14248) );
  MOAI1S U17209 ( .A1(n15698), .A2(n31054), .B1(n15751), .B2(img[1825]), .O(
        n14246) );
  MOAI1S U17210 ( .A1(n15780), .A2(n31096), .B1(n15568), .B2(img[801]), .O(
        n14245) );
  NR2 U17211 ( .I1(n14246), .I2(n14245), .O(n14247) );
  ND3 U17212 ( .I1(n14249), .I2(n14248), .I3(n14247), .O(n16939) );
  ND2S U17213 ( .I1(n16939), .I2(n20620), .O(n14252) );
  ND3 U17214 ( .I1(n14254), .I2(n14253), .I3(n14252), .O(n14255) );
  NR2T U17215 ( .I1(n14256), .I2(n14255), .O(n19554) );
  ND2 U17216 ( .I1(n14257), .I2(n23794), .O(n14258) );
  INV1S U17217 ( .I(n18134), .O(n22927) );
  MOAI1 U17218 ( .A1(n16933), .A2(n15448), .B1(n16932), .B2(n20439), .O(n14265) );
  MOAI1 U17219 ( .A1(n16935), .A2(n13945), .B1(n16934), .B2(n17938), .O(n14264) );
  INV3 U17220 ( .I(n17397), .O(n20124) );
  AOI22S U17221 ( .A1(n16939), .A2(n20124), .B1(n13846), .B2(n16938), .O(
        n14261) );
  BUF1 U17222 ( .I(n17418), .O(n17931) );
  ND2S U17223 ( .I1(n16940), .I2(n17931), .O(n14260) );
  OAI112HS U17224 ( .C1(n14262), .C2(n13766), .A1(n14261), .B1(n14260), .O(
        n14263) );
  NR3H U17225 ( .I1(n14265), .I2(n14264), .I3(n14263), .O(n14285) );
  BUF1 U17226 ( .I(n16059), .O(n17656) );
  AOI22S U17227 ( .A1(n15653), .A2(img[897]), .B1(n15660), .B2(img[129]), .O(
        n14270) );
  AOI22S U17228 ( .A1(n13896), .A2(img[385]), .B1(n15537), .B2(img[257]), .O(
        n14269) );
  AOI22S U17229 ( .A1(n13787), .A2(img[1153]), .B1(n13783), .B2(img[1281]), 
        .O(n14268) );
  AOI22S U17230 ( .A1(n17816), .A2(img[1]), .B1(n15506), .B2(img[513]), .O(
        n14267) );
  AN4S U17231 ( .I1(n14270), .I2(n14269), .I3(n14268), .I4(n14267), .O(n14277)
         );
  MOAI1S U17232 ( .A1(n13850), .A2(n31065), .B1(n15080), .B2(img[1921]), .O(
        n14272) );
  MOAI1S U17233 ( .A1(n15765), .A2(n31053), .B1(n13837), .B2(img[641]), .O(
        n14271) );
  NR2 U17234 ( .I1(n14272), .I2(n14271), .O(n14276) );
  MOAI1S U17235 ( .A1(n15698), .A2(n31061), .B1(n15751), .B2(img[1793]), .O(
        n14274) );
  MOAI1S U17236 ( .A1(n15780), .A2(n31033), .B1(n13885), .B2(img[769]), .O(
        n14273) );
  NR2 U17237 ( .I1(n14274), .I2(n14273), .O(n14275) );
  ND3 U17238 ( .I1(n14277), .I2(n14276), .I3(n14275), .O(n16953) );
  MOAI1 U17239 ( .A1(n16951), .A2(n17656), .B1(n16953), .B2(n13847), .O(n14280) );
  ND2P U17240 ( .I1(n23834), .I2(n14278), .O(n17658) );
  MOAI1 U17241 ( .A1(n16954), .A2(n17658), .B1(n16956), .B2(n13839), .O(n14279) );
  NR2 U17242 ( .I1(n14280), .I2(n14279), .O(n14284) );
  MOAI1 U17243 ( .A1(n16948), .A2(n16468), .B1(n16947), .B2(n20969), .O(n14281) );
  NR2 U17244 ( .I1(n14282), .I2(n14281), .O(n14283) );
  ND3P U17245 ( .I1(n14285), .I2(n14284), .I3(n14283), .O(n14286) );
  MOAI1HP U17246 ( .A1(n19554), .A2(n20969), .B1(n22927), .B2(n13887), .O(
        n21333) );
  INV1S U17247 ( .I(n21333), .O(n15886) );
  NR2 U17248 ( .I1(n21728), .I2(n15886), .O(n15839) );
  INV1S U17249 ( .I(template_store[43]), .O(n15868) );
  MOAI1S U17250 ( .A1(n19648), .A2(n30750), .B1(n19642), .B2(img[154]), .O(
        n14287) );
  AOI22S U17251 ( .A1(n15800), .A2(img[1178]), .B1(n15315), .B2(img[1306]), 
        .O(n14290) );
  AOI22S U17252 ( .A1(n18819), .A2(img[26]), .B1(n15506), .B2(img[538]), .O(
        n14289) );
  AOI22S U17253 ( .A1(n13865), .A2(img[1818]), .B1(n13874), .B2(img[1562]), 
        .O(n14296) );
  MOAI1S U17254 ( .A1(n13850), .A2(n30737), .B1(n22928), .B2(img[1946]), .O(
        n14293) );
  MOAI1S U17255 ( .A1(n14914), .A2(n30677), .B1(n13797), .B2(img[666]), .O(
        n14292) );
  NR2 U17256 ( .I1(n14293), .I2(n14292), .O(n14295) );
  AOI22S U17257 ( .A1(n13885), .A2(img[794]), .B1(n17862), .B2(img[1434]), .O(
        n14294) );
  ND3S U17258 ( .I1(n14296), .I2(n14295), .I3(n14294), .O(n14297) );
  NR2 U17259 ( .I1(n14298), .I2(n14297), .O(n17398) );
  INV1 U17260 ( .I(n14896), .O(n15721) );
  AOI22S U17261 ( .A1(n13882), .A2(img[474]), .B1(n17088), .B2(img[1370]), .O(
        n14302) );
  ND2S U17262 ( .I1(n13885), .I2(img[858]), .O(n14301) );
  ND2S U17263 ( .I1(n15786), .I2(img[346]), .O(n14300) );
  AOI22S U17264 ( .A1(n17515), .A2(img[90]), .B1(n15773), .B2(img[218]), .O(
        n14304) );
  ND2S U17265 ( .I1(n15800), .I2(img[1242]), .O(n14303) );
  OAI112HS U17266 ( .C1(n15698), .C2(n30684), .A1(n14304), .B1(n14303), .O(
        n14305) );
  MOAI1S U17267 ( .A1(n15765), .A2(n30676), .B1(n13797), .B2(img[730]), .O(
        n14308) );
  MOAI1S U17268 ( .A1(n19648), .A2(n30744), .B1(n15657), .B2(img[602]), .O(
        n14307) );
  NR2 U17269 ( .I1(n14308), .I2(n14307), .O(n14312) );
  MOAI1S U17270 ( .A1(n13850), .A2(n30740), .B1(n15080), .B2(img[2010]), .O(
        n14310) );
  NR2 U17271 ( .I1(n14310), .I2(n14309), .O(n14311) );
  ND3 U17272 ( .I1(n14313), .I2(n14312), .I3(n14311), .O(n17396) );
  BUF1 U17273 ( .I(n17418), .O(n20406) );
  MOAI1 U17274 ( .A1(n17398), .A2(n13766), .B1(n17396), .B2(n20406), .O(n14386) );
  MOAI1S U17275 ( .A1(n15674), .A2(n30701), .B1(n15800), .B2(img[1202]), .O(
        n14314) );
  NR2 U17276 ( .I1(n14315), .I2(n14314), .O(n14318) );
  AOI22S U17277 ( .A1(n15537), .A2(img[306]), .B1(n13853), .B2(img[1330]), .O(
        n14317) );
  AOI22S U17278 ( .A1(n13893), .A2(img[946]), .B1(n15506), .B2(img[562]), .O(
        n14316) );
  ND3S U17279 ( .I1(n14318), .I2(n14317), .I3(n14316), .O(n14325) );
  AOI22S U17280 ( .A1(n22928), .A2(img[1970]), .B1(n18148), .B2(img[1074]), 
        .O(n14323) );
  MOAI1S U17281 ( .A1(n15698), .A2(n30575), .B1(n13896), .B2(img[434]), .O(
        n14320) );
  INV1 U17282 ( .I(n19642), .O(n15378) );
  MOAI1S U17283 ( .A1(n15378), .A2(n30705), .B1(n15568), .B2(img[818]), .O(
        n14319) );
  NR2 U17284 ( .I1(n14320), .I2(n14319), .O(n14322) );
  AOI22S U17285 ( .A1(n13898), .A2(img[690]), .B1(n15652), .B2(img[1714]), .O(
        n14321) );
  ND3S U17286 ( .I1(n14323), .I2(n14322), .I3(n14321), .O(n14324) );
  NR2P U17287 ( .I1(n14325), .I2(n14324), .O(n17400) );
  AOI22S U17288 ( .A1(n16048), .A2(img[938]), .B1(n13852), .B2(img[1322]), .O(
        n14329) );
  AOI22S U17289 ( .A1(n22928), .A2(img[1962]), .B1(n15751), .B2(img[1834]), 
        .O(n14328) );
  AOI22S U17290 ( .A1(n15537), .A2(img[298]), .B1(n15773), .B2(img[170]), .O(
        n14327) );
  AOI22S U17291 ( .A1(n13803), .A2(img[42]), .B1(n15800), .B2(img[1194]), .O(
        n14326) );
  AN4S U17292 ( .I1(n14329), .I2(n14328), .I3(n14327), .I4(n14326), .O(n14336)
         );
  MOAI1S U17293 ( .A1(n15765), .A2(n30563), .B1(n13837), .B2(img[682]), .O(
        n14331) );
  MOAI1S U17294 ( .A1(n15277), .A2(n30615), .B1(n13825), .B2(img[554]), .O(
        n14330) );
  NR2 U17295 ( .I1(n14331), .I2(n14330), .O(n14335) );
  MOAI1S U17296 ( .A1(n15780), .A2(n30613), .B1(n13879), .B2(img[426]), .O(
        n14333) );
  OAI22S U17297 ( .A1(n13850), .A2(n30620), .B1(n15698), .B2(n30571), .O(
        n14332) );
  NR2 U17298 ( .I1(n14333), .I2(n14332), .O(n14334) );
  ND3 U17299 ( .I1(n14336), .I2(n14335), .I3(n14334), .O(n17399) );
  MOAI1 U17300 ( .A1(n17400), .A2(n15142), .B1(n17399), .B2(n17875), .O(n14385) );
  MOAI1S U17301 ( .A1(n19648), .A2(n30743), .B1(n19642), .B2(img[162]), .O(
        n14337) );
  NR2 U17302 ( .I1(n14338), .I2(n14337), .O(n14341) );
  AOI22S U17303 ( .A1(n13787), .A2(img[1186]), .B1(n13853), .B2(img[1314]), 
        .O(n14340) );
  AOI22S U17304 ( .A1(n13803), .A2(img[34]), .B1(n15506), .B2(img[546]), .O(
        n14339) );
  ND3 U17305 ( .I1(n14341), .I2(n14340), .I3(n14339), .O(n14348) );
  AOI22S U17306 ( .A1(n13865), .A2(img[1826]), .B1(n15630), .B2(img[1570]), 
        .O(n14346) );
  MOAI1S U17307 ( .A1(n15765), .A2(n30675), .B1(n13837), .B2(img[674]), .O(
        n14342) );
  NR2 U17308 ( .I1(n14343), .I2(n14342), .O(n14345) );
  AOI22S U17309 ( .A1(n19376), .A2(img[802]), .B1(n13845), .B2(img[1442]), .O(
        n14344) );
  ND3S U17310 ( .I1(n14346), .I2(n14345), .I3(n14344), .O(n14347) );
  NR2P U17311 ( .I1(n14348), .I2(n14347), .O(n17405) );
  AOI22S U17312 ( .A1(n13893), .A2(img[898]), .B1(n15773), .B2(img[130]), .O(
        n14352) );
  AOI22S U17313 ( .A1(n13879), .A2(img[386]), .B1(n17578), .B2(img[258]), .O(
        n14351) );
  AOI22S U17314 ( .A1(n15800), .A2(img[1154]), .B1(n13853), .B2(img[1282]), 
        .O(n14350) );
  AOI22S U17315 ( .A1(n13833), .A2(img[2]), .B1(n15506), .B2(img[514]), .O(
        n14349) );
  AN4S U17316 ( .I1(n14352), .I2(n14351), .I3(n14350), .I4(n14349), .O(n14359)
         );
  MOAI1S U17317 ( .A1(n13850), .A2(n30693), .B1(n15080), .B2(img[1922]), .O(
        n14354) );
  MOAI1S U17318 ( .A1(n15765), .A2(n30681), .B1(n13797), .B2(img[642]), .O(
        n14353) );
  NR2 U17319 ( .I1(n14354), .I2(n14353), .O(n14358) );
  MOAI1S U17320 ( .A1(n15698), .A2(n30689), .B1(n15751), .B2(img[1794]), .O(
        n14356) );
  MOAI1S U17321 ( .A1(n15780), .A2(n30662), .B1(n15568), .B2(img[770]), .O(
        n14355) );
  NR2 U17322 ( .I1(n14356), .I2(n14355), .O(n14357) );
  ND3 U17323 ( .I1(n14359), .I2(n14358), .I3(n14357), .O(n17404) );
  INV2 U17324 ( .I(n14259), .O(n21062) );
  AOI22S U17325 ( .A1(n15653), .A2(img[994]), .B1(n15773), .B2(img[226]), .O(
        n14363) );
  AOI22S U17326 ( .A1(n13882), .A2(img[482]), .B1(n19710), .B2(img[354]), .O(
        n14362) );
  AOI22S U17327 ( .A1(n15800), .A2(img[1250]), .B1(n13853), .B2(img[1378]), 
        .O(n14361) );
  AOI22S U17328 ( .A1(n17793), .A2(img[98]), .B1(n13876), .B2(img[610]), .O(
        n14360) );
  MOAI1S U17329 ( .A1(n13850), .A2(n30738), .B1(n15080), .B2(img[2018]), .O(
        n14365) );
  MOAI1S U17330 ( .A1(n15765), .A2(n30678), .B1(n13898), .B2(img[738]), .O(
        n14364) );
  NR2 U17331 ( .I1(n14365), .I2(n14364), .O(n14369) );
  MOAI1S U17332 ( .A1(n15698), .A2(n30686), .B1(n15751), .B2(img[1890]), .O(
        n14367) );
  MOAI1S U17333 ( .A1(n15780), .A2(n30731), .B1(n15568), .B2(img[866]), .O(
        n14366) );
  NR2 U17334 ( .I1(n14367), .I2(n14366), .O(n14368) );
  ND3 U17335 ( .I1(n14370), .I2(n14369), .I3(n14368), .O(n17403) );
  AOI22S U17336 ( .A1(n13893), .A2(img[962]), .B1(n15773), .B2(img[194]), .O(
        n14374) );
  AOI22S U17337 ( .A1(n13882), .A2(img[450]), .B1(n13829), .B2(img[322]), .O(
        n14373) );
  AOI22S U17338 ( .A1(n15800), .A2(img[1218]), .B1(n15315), .B2(img[1346]), 
        .O(n14372) );
  AOI22S U17339 ( .A1(n17886), .A2(img[66]), .B1(n13876), .B2(img[578]), .O(
        n14371) );
  MOAI1S U17340 ( .A1(n13850), .A2(n30692), .B1(n15080), .B2(img[1986]), .O(
        n14376) );
  MOAI1S U17341 ( .A1(n15765), .A2(n30680), .B1(n13837), .B2(img[706]), .O(
        n14375) );
  NR2 U17342 ( .I1(n14376), .I2(n14375), .O(n14380) );
  MOAI1S U17343 ( .A1(n15698), .A2(n30688), .B1(n15751), .B2(img[1858]), .O(
        n14378) );
  MOAI1S U17344 ( .A1(n15780), .A2(n30661), .B1(n15568), .B2(img[834]), .O(
        n14377) );
  NR2 U17345 ( .I1(n14378), .I2(n14377), .O(n14379) );
  ND3 U17346 ( .I1(n14381), .I2(n14380), .I3(n14379), .O(n17407) );
  BUF1 U17347 ( .I(n18040), .O(n20150) );
  ND2S U17348 ( .I1(n17407), .I2(n20150), .O(n14382) );
  OAI112HS U17349 ( .C1(n17405), .C2(n17397), .A1(n14383), .B1(n14382), .O(
        n14384) );
  NR3HP U17350 ( .I1(n14386), .I2(n14385), .I3(n14384), .O(n14488) );
  MOAI1S U17351 ( .A1(n13850), .A2(n30581), .B1(n15080), .B2(img[2034]), .O(
        n14388) );
  MOAI1S U17352 ( .A1(n15698), .A2(n30577), .B1(n13896), .B2(img[498]), .O(
        n14387) );
  NR2 U17353 ( .I1(n14388), .I2(n14387), .O(n14391) );
  MAOI1S U17354 ( .A1(n13898), .A2(img[754]), .B1(n30569), .B2(n15765), .O(
        n14390) );
  INV1S U17355 ( .I(n16758), .O(n16075) );
  AOI22S U17356 ( .A1(n16075), .A2(img[1906]), .B1(n13885), .B2(img[882]), .O(
        n14389) );
  ND3 U17357 ( .I1(n14391), .I2(n14390), .I3(n14389), .O(n14399) );
  MOAI1S U17358 ( .A1(n15780), .A2(n30550), .B1(n19642), .B2(img[242]), .O(
        n14394) );
  NR2 U17359 ( .I1(n14394), .I2(n14393), .O(n14397) );
  AOI22S U17360 ( .A1(n13880), .A2(img[1010]), .B1(n13876), .B2(img[626]), .O(
        n14396) );
  AOI22S U17361 ( .A1(n18996), .A2(img[114]), .B1(n15800), .B2(img[1266]), .O(
        n14395) );
  MOAI1S U17362 ( .A1(n15780), .A2(n30663), .B1(n13879), .B2(img[506]), .O(
        n14405) );
  AOI22S U17363 ( .A1(n22928), .A2(img[2042]), .B1(n15800), .B2(img[1274]), 
        .O(n14402) );
  ND2S U17364 ( .I1(n15657), .I2(img[634]), .O(n14401) );
  ND2S U17365 ( .I1(n17088), .I2(img[1402]), .O(n14400) );
  NR3 U17366 ( .I1(n14405), .I2(n14404), .I3(n14403), .O(n14412) );
  MOAI1S U17367 ( .A1(n18109), .A2(n30674), .B1(n15568), .B2(img[890]), .O(
        n14407) );
  OAI22S U17368 ( .A1(n13850), .A2(n30694), .B1(n15698), .B2(n30690), .O(
        n14406) );
  NR2 U17369 ( .I1(n14407), .I2(n14406), .O(n14411) );
  MOAI1S U17370 ( .A1(n19648), .A2(n30698), .B1(n19290), .B2(img[122]), .O(
        n14409) );
  MOAI1S U17371 ( .A1(n15765), .A2(n30682), .B1(n13797), .B2(img[762]), .O(
        n14408) );
  NR2 U17372 ( .I1(n14409), .I2(n14408), .O(n14410) );
  ND3 U17373 ( .I1(n14412), .I2(n14411), .I3(n14410), .O(n17411) );
  MOAI1 U17374 ( .A1(n17412), .A2(n13947), .B1(n17411), .B2(n20969), .O(n14437) );
  MOAI1S U17375 ( .A1(n15698), .A2(n30576), .B1(n15080), .B2(img[1994]), .O(
        n14414) );
  MOAI1S U17376 ( .A1(n15674), .A2(n30702), .B1(n15657), .B2(img[586]), .O(
        n14413) );
  NR2 U17377 ( .I1(n14414), .I2(n14413), .O(n14417) );
  AOI22S U17378 ( .A1(n13880), .A2(img[970]), .B1(n15773), .B2(img[202]), .O(
        n14416) );
  AOI22S U17379 ( .A1(n13787), .A2(img[1226]), .B1(n13824), .B2(img[1354]), 
        .O(n14415) );
  ND3S U17380 ( .I1(n14417), .I2(n14416), .I3(n14415), .O(n14424) );
  MOAI1S U17381 ( .A1(n13850), .A2(n30580), .B1(n15786), .B2(img[330]), .O(
        n14419) );
  MOAI1S U17382 ( .A1(n15765), .A2(n30568), .B1(n13837), .B2(img[714]), .O(
        n14418) );
  NR2 U17383 ( .I1(n14419), .I2(n14418), .O(n14422) );
  AOI22S U17384 ( .A1(n13786), .A2(img[1866]), .B1(n19641), .B2(img[842]), .O(
        n14421) );
  INV3 U17385 ( .I(n14739), .O(n15780) );
  ND3 U17386 ( .I1(n14422), .I2(n14421), .I3(n14420), .O(n14423) );
  AOI22S U17387 ( .A1(n13893), .A2(img[1002]), .B1(n15773), .B2(img[234]), .O(
        n14428) );
  AOI22S U17388 ( .A1(n18262), .A2(img[490]), .B1(n19018), .B2(img[362]), .O(
        n14427) );
  AOI22S U17389 ( .A1(n18922), .A2(img[1258]), .B1(n15315), .B2(img[1386]), 
        .O(n14426) );
  AOI22S U17390 ( .A1(n18996), .A2(img[106]), .B1(n15506), .B2(img[618]), .O(
        n14425) );
  MOAI1S U17391 ( .A1(n13850), .A2(n30619), .B1(n15080), .B2(img[2026]), .O(
        n14430) );
  MOAI1S U17392 ( .A1(n15765), .A2(n30566), .B1(n13797), .B2(img[746]), .O(
        n14429) );
  NR2 U17393 ( .I1(n14430), .I2(n14429), .O(n14434) );
  MOAI1S U17394 ( .A1(n15698), .A2(n30574), .B1(n15751), .B2(img[1898]), .O(
        n14432) );
  MOAI1S U17395 ( .A1(n15780), .A2(n30612), .B1(n15568), .B2(img[874]), .O(
        n14431) );
  NR2 U17396 ( .I1(n14432), .I2(n14431), .O(n14433) );
  NR2 U17397 ( .I1(n14437), .I2(n14436), .O(n14487) );
  AOI22S U17398 ( .A1(n13845), .A2(img[1426]), .B1(n13874), .B2(img[1554]), 
        .O(n14442) );
  MOAI1S U17399 ( .A1(n13850), .A2(n30618), .B1(n15080), .B2(img[1938]), .O(
        n14439) );
  MOAI1S U17400 ( .A1(n15765), .A2(n30565), .B1(n13837), .B2(img[658]), .O(
        n14438) );
  NR2 U17401 ( .I1(n14439), .I2(n14438), .O(n14441) );
  AOI22S U17402 ( .A1(n15660), .A2(img[146]), .B1(n19376), .B2(img[786]), .O(
        n14440) );
  MOAI1S U17403 ( .A1(n19648), .A2(n30631), .B1(n13876), .B2(img[530]), .O(
        n14444) );
  MOAI1S U17404 ( .A1(n14896), .A2(n30635), .B1(n15800), .B2(img[1170]), .O(
        n14443) );
  NR2 U17405 ( .I1(n14444), .I2(n14443), .O(n14447) );
  AOI22S U17406 ( .A1(n15537), .A2(img[274]), .B1(n13801), .B2(img[18]), .O(
        n14446) );
  AOI22S U17407 ( .A1(n19036), .A2(img[1810]), .B1(n15315), .B2(img[1298]), 
        .O(n14445) );
  ND3S U17408 ( .I1(n14447), .I2(n14446), .I3(n14445), .O(n14448) );
  AOI22S U17409 ( .A1(n13893), .A2(img[978]), .B1(n15773), .B2(img[210]), .O(
        n14453) );
  AOI22S U17410 ( .A1(n13896), .A2(img[466]), .B1(n17534), .B2(img[338]), .O(
        n14452) );
  AOI22S U17411 ( .A1(n15800), .A2(img[1234]), .B1(n17088), .B2(img[1362]), 
        .O(n14451) );
  AOI22S U17412 ( .A1(n18773), .A2(img[82]), .B1(n15506), .B2(img[594]), .O(
        n14450) );
  MOAI1S U17413 ( .A1(n13850), .A2(n30621), .B1(n15080), .B2(img[2002]), .O(
        n14455) );
  MOAI1S U17414 ( .A1(n15765), .A2(n30564), .B1(n13837), .B2(img[722]), .O(
        n14454) );
  NR2 U17415 ( .I1(n14455), .I2(n14454), .O(n14459) );
  MOAI1S U17416 ( .A1(n15698), .A2(n30572), .B1(n15751), .B2(img[1874]), .O(
        n14457) );
  MOAI1S U17417 ( .A1(n15780), .A2(n30614), .B1(n15568), .B2(img[850]), .O(
        n14456) );
  NR2 U17418 ( .I1(n14457), .I2(n14456), .O(n14458) );
  ND3 U17419 ( .I1(n14460), .I2(n14459), .I3(n14458), .O(n17419) );
  MOAI1 U17420 ( .A1(n17417), .A2(n17656), .B1(n17419), .B2(n17938), .O(n14485) );
  MOAI1S U17421 ( .A1(n13894), .A2(n30770), .B1(n15786), .B2(img[314]), .O(
        n14462) );
  MOAI1S U17422 ( .A1(n19648), .A2(n30764), .B1(n19642), .B2(img[186]), .O(
        n14461) );
  AOI22S U17423 ( .A1(n18838), .A2(img[1210]), .B1(n13853), .B2(img[1338]), 
        .O(n14464) );
  AOI22S U17424 ( .A1(n19411), .A2(img[58]), .B1(n20102), .B2(img[570]), .O(
        n14463) );
  ND3 U17425 ( .I1(n14465), .I2(n14464), .I3(n14463), .O(n14472) );
  AOI22S U17426 ( .A1(n19036), .A2(img[1850]), .B1(n19193), .B2(img[1594]), 
        .O(n14470) );
  MOAI1S U17427 ( .A1(n13850), .A2(n30691), .B1(n15080), .B2(img[1978]), .O(
        n14467) );
  MOAI1S U17428 ( .A1(n15765), .A2(n30679), .B1(n13837), .B2(img[698]), .O(
        n14466) );
  NR2 U17429 ( .I1(n14467), .I2(n14466), .O(n14469) );
  AOI22S U17430 ( .A1(n13875), .A2(img[826]), .B1(n13845), .B2(img[1466]), .O(
        n14468) );
  ND3S U17431 ( .I1(n14470), .I2(n14469), .I3(n14468), .O(n14471) );
  AOI22S U17432 ( .A1(n16048), .A2(img[906]), .B1(n15773), .B2(img[138]), .O(
        n14476) );
  AOI22S U17433 ( .A1(n13896), .A2(img[394]), .B1(n18796), .B2(img[266]), .O(
        n14475) );
  AOI22S U17434 ( .A1(n18922), .A2(img[1162]), .B1(n15315), .B2(img[1290]), 
        .O(n14474) );
  AOI22S U17435 ( .A1(n17886), .A2(img[10]), .B1(n13785), .B2(img[522]), .O(
        n14473) );
  AN4S U17436 ( .I1(n14476), .I2(n14475), .I3(n14474), .I4(n14473), .O(n14483)
         );
  MOAI1S U17437 ( .A1(n13850), .A2(n30582), .B1(n15080), .B2(img[1930]), .O(
        n14478) );
  MOAI1S U17438 ( .A1(n15765), .A2(n30570), .B1(n13837), .B2(img[650]), .O(
        n14477) );
  NR2 U17439 ( .I1(n14478), .I2(n14477), .O(n14482) );
  MOAI1S U17440 ( .A1(n15698), .A2(n30578), .B1(n15751), .B2(img[1802]), .O(
        n14480) );
  MOAI1S U17441 ( .A1(n15780), .A2(n30551), .B1(n15568), .B2(img[778]), .O(
        n14479) );
  NR2 U17442 ( .I1(n14480), .I2(n14479), .O(n14481) );
  ND3 U17443 ( .I1(n14483), .I2(n14482), .I3(n14481), .O(n17422) );
  MOAI1 U17444 ( .A1(n17421), .A2(n17658), .B1(n17422), .B2(n13830), .O(n14484) );
  ND3HT U17445 ( .I1(n14488), .I2(n14487), .I3(n14486), .O(n21225) );
  INV1S U17446 ( .I(n17411), .O(n14489) );
  MOAI1S U17447 ( .A1(n14489), .A2(n13947), .B1(n17396), .B2(n17938), .O(
        n14491) );
  INV2 U17448 ( .I(n17397), .O(n20613) );
  NR2 U17449 ( .I1(n14491), .I2(n14490), .O(n14494) );
  AOI22S U17450 ( .A1(n17413), .A2(n21062), .B1(n20263), .B2(n17419), .O(
        n14492) );
  ND3S U17451 ( .I1(n14494), .I2(n14493), .I3(n14492), .O(n14502) );
  OAI22S U17452 ( .A1(n17405), .A2(n13766), .B1(n17414), .B2(n20421), .O(
        n14495) );
  NR2 U17453 ( .I1(n14496), .I2(n14495), .O(n14500) );
  INV1S U17454 ( .I(n17398), .O(n14497) );
  AOI22S U17455 ( .A1(n13843), .A2(n17407), .B1(n14497), .B2(n17762), .O(
        n14499) );
  ND2S U17456 ( .I1(n17422), .I2(n13847), .O(n14498) );
  ND3 U17457 ( .I1(n14500), .I2(n14499), .I3(n14498), .O(n14501) );
  NR2 U17458 ( .I1(n14502), .I2(n14501), .O(n14503) );
  INV1S U17459 ( .I(n19534), .O(n14504) );
  OAI12H U17460 ( .B1(n13818), .B2(n18134), .A1(n14504), .O(n20436) );
  INV2 U17461 ( .I(n20436), .O(n15867) );
  NR2 U17462 ( .I1(n15868), .I2(n15867), .O(n15372) );
  MOAI1S U17463 ( .A1(n13850), .A2(n31548), .B1(n15080), .B2(img[2040]), .O(
        n14507) );
  MOAI1S U17464 ( .A1(n15765), .A2(n31536), .B1(n13797), .B2(img[760]), .O(
        n14506) );
  NR2 U17465 ( .I1(n14507), .I2(n14506), .O(n14510) );
  AOI22S U17466 ( .A1(n15537), .A2(img[376]), .B1(n13885), .B2(img[888]), .O(
        n14508) );
  ND3S U17467 ( .I1(n14510), .I2(n14509), .I3(n14508), .O(n14517) );
  MOAI1S U17468 ( .A1(n15668), .A2(n31512), .B1(n15800), .B2(img[1272]), .O(
        n14512) );
  MOAI1S U17469 ( .A1(n19648), .A2(n31563), .B1(n15657), .B2(img[632]), .O(
        n14511) );
  NR2 U17470 ( .I1(n14512), .I2(n14511), .O(n14515) );
  AOI22S U17471 ( .A1(n19411), .A2(img[120]), .B1(n13783), .B2(img[1400]), .O(
        n14514) );
  AOI22S U17472 ( .A1(n13896), .A2(img[504]), .B1(n15660), .B2(img[248]), .O(
        n14513) );
  ND3S U17473 ( .I1(n14515), .I2(n14514), .I3(n14513), .O(n14516) );
  NR2 U17474 ( .I1(n14517), .I2(n14516), .O(n14716) );
  AOI22S U17475 ( .A1(n18718), .A2(img[1008]), .B1(n15660), .B2(img[240]), .O(
        n14521) );
  AOI22S U17476 ( .A1(n13896), .A2(img[496]), .B1(n15537), .B2(img[368]), .O(
        n14520) );
  AOI22S U17477 ( .A1(n15800), .A2(img[1264]), .B1(n14392), .B2(img[1392]), 
        .O(n14519) );
  AOI22S U17478 ( .A1(n13803), .A2(img[112]), .B1(n15506), .B2(img[624]), .O(
        n14518) );
  AN4S U17479 ( .I1(n14521), .I2(n14520), .I3(n14519), .I4(n14518), .O(n14528)
         );
  MOAI1S U17480 ( .A1(n13850), .A2(n31665), .B1(n15080), .B2(img[2032]), .O(
        n14523) );
  MOAI1S U17481 ( .A1(n15765), .A2(n31611), .B1(n13797), .B2(img[752]), .O(
        n14522) );
  NR2 U17482 ( .I1(n14523), .I2(n14522), .O(n14527) );
  MOAI1S U17483 ( .A1(n15698), .A2(n31619), .B1(n15809), .B2(img[1904]), .O(
        n14525) );
  MOAI1S U17484 ( .A1(n15780), .A2(n31658), .B1(n13885), .B2(img[880]), .O(
        n14524) );
  NR2 U17485 ( .I1(n14525), .I2(n14524), .O(n14526) );
  ND3 U17486 ( .I1(n14528), .I2(n14527), .I3(n14526), .O(n17166) );
  MOAI1 U17487 ( .A1(n14716), .A2(n13844), .B1(n17166), .B2(n13846), .O(n14603) );
  MOAI1S U17488 ( .A1(n13850), .A2(n31626), .B1(n15080), .B2(img[1936]), .O(
        n14530) );
  MOAI1S U17489 ( .A1(n15780), .A2(n31595), .B1(n15809), .B2(img[1808]), .O(
        n14529) );
  NR2 U17490 ( .I1(n14530), .I2(n14529), .O(n14533) );
  AOI22S U17491 ( .A1(n13898), .A2(img[656]), .B1(n15652), .B2(img[1680]), .O(
        n14532) );
  AOI22S U17492 ( .A1(n15537), .A2(img[272]), .B1(n13884), .B2(img[784]), .O(
        n14531) );
  ND3 U17493 ( .I1(n14533), .I2(n14532), .I3(n14531), .O(n14540) );
  MOAI1S U17494 ( .A1(n15698), .A2(n31622), .B1(n15653), .B2(img[912]), .O(
        n14535) );
  MOAI1S U17495 ( .A1(n15674), .A2(n31575), .B1(n15657), .B2(img[528]), .O(
        n14534) );
  NR2 U17496 ( .I1(n14535), .I2(n14534), .O(n14538) );
  AOI22S U17497 ( .A1(n13896), .A2(img[400]), .B1(n15660), .B2(img[144]), .O(
        n14537) );
  AOI22S U17498 ( .A1(n15800), .A2(img[1168]), .B1(n18729), .B2(img[1296]), 
        .O(n14536) );
  ND3S U17499 ( .I1(n14538), .I2(n14537), .I3(n14536), .O(n14539) );
  NR2 U17500 ( .I1(n14540), .I2(n14539), .O(n14709) );
  MOAI1S U17501 ( .A1(n13850), .A2(n31550), .B1(n15080), .B2(img[1984]), .O(
        n14545) );
  MOAI1S U17502 ( .A1(n15765), .A2(n31538), .B1(n13797), .B2(img[704]), .O(
        n14544) );
  AOI22S U17503 ( .A1(n15691), .A2(img[448]), .B1(n15537), .B2(img[320]), .O(
        n14542) );
  ND2S U17504 ( .I1(n13884), .I2(img[832]), .O(n14541) );
  OAI112HS U17505 ( .C1(n15698), .C2(n31546), .A1(n14542), .B1(n14541), .O(
        n14543) );
  NR3 U17506 ( .I1(n14545), .I2(n14544), .I3(n14543), .O(n14552) );
  MOAI1S U17507 ( .A1(n19648), .A2(n31522), .B1(n19642), .B2(img[192]), .O(
        n14547) );
  MOAI1S U17508 ( .A1(n13789), .A2(n31520), .B1(n13841), .B2(img[64]), .O(
        n14546) );
  NR2 U17509 ( .I1(n14547), .I2(n14546), .O(n14551) );
  MOAI1S U17510 ( .A1(n18109), .A2(n31508), .B1(n15800), .B2(img[1216]), .O(
        n14549) );
  MOAI1S U17511 ( .A1(n15780), .A2(n31514), .B1(n15657), .B2(img[576]), .O(
        n14548) );
  NR2 U17512 ( .I1(n14549), .I2(n14548), .O(n14550) );
  ND3 U17513 ( .I1(n14552), .I2(n14551), .I3(n14550), .O(n17160) );
  MOAI1 U17514 ( .A1(n14709), .A2(n17656), .B1(n17160), .B2(n18040), .O(n14602) );
  MOAI1S U17515 ( .A1(n19648), .A2(n31731), .B1(n19642), .B2(img[152]), .O(
        n14553) );
  NR2 U17516 ( .I1(n14554), .I2(n14553), .O(n14558) );
  AOI22S U17517 ( .A1(n15561), .A2(img[1176]), .B1(n13824), .B2(img[1304]), 
        .O(n14557) );
  AOI22S U17518 ( .A1(n18773), .A2(img[24]), .B1(n15657), .B2(img[536]), .O(
        n14556) );
  AOI22S U17519 ( .A1(n19023), .A2(img[1816]), .B1(n15630), .B2(img[1560]), 
        .O(n14563) );
  MOAI1S U17520 ( .A1(n13850), .A2(n31694), .B1(n15080), .B2(img[1944]), .O(
        n14560) );
  MOAI1S U17521 ( .A1(n15765), .A2(n31533), .B1(n13797), .B2(img[664]), .O(
        n14559) );
  NR2 U17522 ( .I1(n14560), .I2(n14559), .O(n14562) );
  AOI22S U17523 ( .A1(n13875), .A2(img[792]), .B1(n13845), .B2(img[1432]), .O(
        n14561) );
  ND3S U17524 ( .I1(n14563), .I2(n14562), .I3(n14561), .O(n14564) );
  AOI22S U17525 ( .A1(n13892), .A2(img[896]), .B1(n15660), .B2(img[128]), .O(
        n14569) );
  AOI22S U17526 ( .A1(n13896), .A2(img[384]), .B1(n15537), .B2(img[256]), .O(
        n14568) );
  AOI22S U17527 ( .A1(n15561), .A2(img[1152]), .B1(n13854), .B2(img[1280]), 
        .O(n14567) );
  AOI22S U17528 ( .A1(n18958), .A2(img[0]), .B1(n15657), .B2(img[512]), .O(
        n14566) );
  AN4S U17529 ( .I1(n14569), .I2(n14568), .I3(n14567), .I4(n14566), .O(n14576)
         );
  MOAI1S U17530 ( .A1(n13850), .A2(n31547), .B1(n15080), .B2(img[1920]), .O(
        n14571) );
  MOAI1S U17531 ( .A1(n15765), .A2(n31535), .B1(n13837), .B2(img[640]), .O(
        n14570) );
  NR2 U17532 ( .I1(n14571), .I2(n14570), .O(n14575) );
  MOAI1S U17533 ( .A1(n15698), .A2(n31543), .B1(n15809), .B2(img[1792]), .O(
        n14573) );
  MOAI1S U17534 ( .A1(n15668), .A2(n31511), .B1(n13885), .B2(img[768]), .O(
        n14572) );
  NR2 U17535 ( .I1(n14573), .I2(n14572), .O(n14574) );
  ND3 U17536 ( .I1(n14576), .I2(n14575), .I3(n14574), .O(n17171) );
  AOI22S U17537 ( .A1(n15653), .A2(img[992]), .B1(n15660), .B2(img[224]), .O(
        n14580) );
  AOI22S U17538 ( .A1(n13879), .A2(img[480]), .B1(n15537), .B2(img[352]), .O(
        n14579) );
  AOI22S U17539 ( .A1(n15561), .A2(img[1248]), .B1(n15315), .B2(img[1376]), 
        .O(n14578) );
  AOI22S U17540 ( .A1(n13803), .A2(img[96]), .B1(n15657), .B2(img[608]), .O(
        n14577) );
  MOAI1S U17541 ( .A1(n13850), .A2(n31695), .B1(n15080), .B2(img[2016]), .O(
        n14582) );
  NR2 U17542 ( .I1(n14582), .I2(n14581), .O(n14586) );
  MOAI1S U17543 ( .A1(n15698), .A2(n31542), .B1(n15809), .B2(img[1888]), .O(
        n14584) );
  NR2 U17544 ( .I1(n14584), .I2(n14583), .O(n14585) );
  AOI22S U17545 ( .A1(n17171), .A2(n13847), .B1(n21062), .B2(n17178), .O(
        n14600) );
  AOI22S U17546 ( .A1(n19403), .A2(img[968]), .B1(n15660), .B2(img[200]), .O(
        n14591) );
  AOI22S U17547 ( .A1(n13896), .A2(img[456]), .B1(n18736), .B2(img[328]), .O(
        n14590) );
  AOI22S U17548 ( .A1(n15561), .A2(img[1224]), .B1(n13854), .B2(img[1352]), 
        .O(n14589) );
  AOI22S U17549 ( .A1(n18958), .A2(img[72]), .B1(n13883), .B2(img[584]), .O(
        n14588) );
  MOAI1S U17550 ( .A1(n13850), .A2(n31664), .B1(n15080), .B2(img[1992]), .O(
        n14593) );
  MOAI1S U17551 ( .A1(n15765), .A2(n31609), .B1(n13837), .B2(img[712]), .O(
        n14592) );
  NR2 U17552 ( .I1(n14593), .I2(n14592), .O(n14597) );
  MOAI1S U17553 ( .A1(n15698), .A2(n31617), .B1(n15809), .B2(img[1864]), .O(
        n14595) );
  MOAI1S U17554 ( .A1(n15780), .A2(n31657), .B1(n13885), .B2(img[840]), .O(
        n14594) );
  NR2 U17555 ( .I1(n14595), .I2(n14594), .O(n14596) );
  ND3 U17556 ( .I1(n14598), .I2(n14597), .I3(n14596), .O(n17173) );
  ND2S U17557 ( .I1(n17173), .I2(n20439), .O(n14599) );
  OAI112HS U17558 ( .C1(n17172), .C2(n13766), .A1(n14600), .B1(n14599), .O(
        n14601) );
  MOAI1S U17559 ( .A1(n19648), .A2(n31716), .B1(n19642), .B2(img[176]), .O(
        n14604) );
  NR2 U17560 ( .I1(n14605), .I2(n14604), .O(n14608) );
  AOI22S U17561 ( .A1(n15561), .A2(img[1200]), .B1(n18824), .B2(img[1328]), 
        .O(n14607) );
  AOI22S U17562 ( .A1(n18773), .A2(img[48]), .B1(n15506), .B2(img[560]), .O(
        n14606) );
  ND3 U17563 ( .I1(n14608), .I2(n14607), .I3(n14606), .O(n14615) );
  AOI22S U17564 ( .A1(n13863), .A2(img[1840]), .B1(n20109), .B2(img[1584]), 
        .O(n14613) );
  MOAI1S U17565 ( .A1(n13850), .A2(n31663), .B1(n15080), .B2(img[1968]), .O(
        n14610) );
  MOAI1S U17566 ( .A1(n15765), .A2(n31608), .B1(n13898), .B2(img[688]), .O(
        n14609) );
  NR2 U17567 ( .I1(n14610), .I2(n14609), .O(n14612) );
  AOI22S U17568 ( .A1(n13884), .A2(img[816]), .B1(n13845), .B2(img[1456]), .O(
        n14611) );
  ND3S U17569 ( .I1(n14613), .I2(n14612), .I3(n14611), .O(n14614) );
  NR2P U17570 ( .I1(n14615), .I2(n14614), .O(n17174) );
  AOI22S U17571 ( .A1(n13896), .A2(img[464]), .B1(n13853), .B2(img[1360]), .O(
        n14618) );
  ND2S U17572 ( .I1(n13892), .I2(img[976]), .O(n14617) );
  ND2S U17573 ( .I1(n15657), .I2(img[592]), .O(n14616) );
  ND3S U17574 ( .I1(n14618), .I2(n14617), .I3(n14616), .O(n14622) );
  AOI22S U17575 ( .A1(n13803), .A2(img[80]), .B1(n15800), .B2(img[1232]), .O(
        n14620) );
  ND2S U17576 ( .I1(n19642), .I2(img[208]), .O(n14619) );
  OAI112HS U17577 ( .C1(n13850), .C2(n31625), .A1(n14620), .B1(n14619), .O(
        n14621) );
  NR2 U17578 ( .I1(n14622), .I2(n14621), .O(n14629) );
  MOAI1S U17579 ( .A1(n15698), .A2(n31621), .B1(n15080), .B2(img[2000]), .O(
        n14624) );
  MOAI1S U17580 ( .A1(n15765), .A2(n31613), .B1(n13898), .B2(img[720]), .O(
        n14623) );
  NR2 U17581 ( .I1(n14624), .I2(n14623), .O(n14628) );
  MOAI1S U17582 ( .A1(n15631), .A2(n31706), .B1(n13885), .B2(img[848]), .O(
        n14625) );
  NR2 U17583 ( .I1(n14626), .I2(n14625), .O(n14627) );
  ND3 U17584 ( .I1(n14629), .I2(n14628), .I3(n14627), .O(n17167) );
  MOAI1 U17585 ( .A1(n17174), .A2(n15142), .B1(n17167), .B2(n17938), .O(n14654) );
  MOAI1S U17586 ( .A1(n15113), .A2(n31527), .B1(n15786), .B2(img[312]), .O(
        n14631) );
  MOAI1S U17587 ( .A1(n19648), .A2(n31521), .B1(n19642), .B2(img[184]), .O(
        n14630) );
  AOI22S U17588 ( .A1(n15561), .A2(img[1208]), .B1(n16799), .B2(img[1336]), 
        .O(n14633) );
  AOI22S U17589 ( .A1(n13803), .A2(img[56]), .B1(n15506), .B2(img[568]), .O(
        n14632) );
  AOI22S U17590 ( .A1(n19036), .A2(img[1848]), .B1(n15630), .B2(img[1592]), 
        .O(n14639) );
  MOAI1S U17591 ( .A1(n13850), .A2(n31549), .B1(n15080), .B2(img[1976]), .O(
        n14636) );
  MOAI1S U17592 ( .A1(n15765), .A2(n31537), .B1(n13837), .B2(img[696]), .O(
        n14635) );
  NR2 U17593 ( .I1(n14636), .I2(n14635), .O(n14638) );
  AOI22S U17594 ( .A1(n16348), .A2(img[824]), .B1(n13845), .B2(img[1464]), .O(
        n14637) );
  ND3S U17595 ( .I1(n14639), .I2(n14638), .I3(n14637), .O(n14640) );
  AOI22S U17596 ( .A1(n15653), .A2(img[928]), .B1(n15800), .B2(img[1184]), .O(
        n14645) );
  AOI22S U17597 ( .A1(n15691), .A2(img[416]), .B1(n15537), .B2(img[288]), .O(
        n14644) );
  AOI22S U17598 ( .A1(n13801), .A2(img[32]), .B1(n13785), .B2(img[544]), .O(
        n14643) );
  AOI22S U17599 ( .A1(n15660), .A2(img[160]), .B1(n13783), .B2(img[1312]), .O(
        n14642) );
  AN4S U17600 ( .I1(n14645), .I2(n14644), .I3(n14643), .I4(n14642), .O(n14652)
         );
  MOAI1S U17601 ( .A1(n15765), .A2(n31531), .B1(n13797), .B2(img[672]), .O(
        n14647) );
  MOAI1S U17602 ( .A1(n13850), .A2(n31696), .B1(n13885), .B2(img[800]), .O(
        n14646) );
  NR2 U17603 ( .I1(n14647), .I2(n14646), .O(n14651) );
  MOAI1S U17604 ( .A1(n15698), .A2(n31539), .B1(n15080), .B2(img[1952]), .O(
        n14649) );
  MOAI1S U17605 ( .A1(n15780), .A2(n31689), .B1(n15809), .B2(img[1824]), .O(
        n14648) );
  NR2 U17606 ( .I1(n14649), .I2(n14648), .O(n14650) );
  ND3 U17607 ( .I1(n14652), .I2(n14651), .I3(n14650), .O(n17180) );
  MOAI1 U17608 ( .A1(n17165), .A2(n17658), .B1(n17180), .B2(n20613), .O(n14653) );
  NR2P U17609 ( .I1(n14654), .I2(n14653), .O(n14704) );
  MOAI1S U17610 ( .A1(n19648), .A2(n31649), .B1(n19642), .B2(img[136]), .O(
        n14655) );
  NR2 U17611 ( .I1(n14656), .I2(n14655), .O(n14659) );
  AOI22S U17612 ( .A1(n15561), .A2(img[1160]), .B1(n13853), .B2(img[1288]), 
        .O(n14658) );
  AOI22S U17613 ( .A1(n13833), .A2(img[8]), .B1(n13785), .B2(img[520]), .O(
        n14657) );
  AOI22S U17614 ( .A1(n13865), .A2(img[1800]), .B1(n15630), .B2(img[1544]), 
        .O(n14664) );
  MOAI1S U17615 ( .A1(n13850), .A2(n31666), .B1(n15080), .B2(img[1928]), .O(
        n14661) );
  MOAI1S U17616 ( .A1(n15765), .A2(n31610), .B1(n13837), .B2(img[648]), .O(
        n14660) );
  NR2 U17617 ( .I1(n14661), .I2(n14660), .O(n14663) );
  AOI22S U17618 ( .A1(n16348), .A2(img[776]), .B1(n13845), .B2(img[1416]), .O(
        n14662) );
  ND3S U17619 ( .I1(n14664), .I2(n14663), .I3(n14662), .O(n14665) );
  AOI22S U17620 ( .A1(n13893), .A2(img[984]), .B1(n15660), .B2(img[216]), .O(
        n14670) );
  AOI22S U17621 ( .A1(n15691), .A2(img[472]), .B1(n15537), .B2(img[344]), .O(
        n14669) );
  AOI22S U17622 ( .A1(n15561), .A2(img[1240]), .B1(n13853), .B2(img[1368]), 
        .O(n14668) );
  AOI22S U17623 ( .A1(n17816), .A2(img[88]), .B1(n13876), .B2(img[600]), .O(
        n14667) );
  AN4S U17624 ( .I1(n14670), .I2(n14669), .I3(n14668), .I4(n14667), .O(n14677)
         );
  MOAI1S U17625 ( .A1(n13850), .A2(n31697), .B1(n15080), .B2(img[2008]), .O(
        n14672) );
  MOAI1S U17626 ( .A1(n15765), .A2(n31532), .B1(n13837), .B2(img[728]), .O(
        n14671) );
  NR2 U17627 ( .I1(n14672), .I2(n14671), .O(n14676) );
  MOAI1S U17628 ( .A1(n15698), .A2(n31540), .B1(n15809), .B2(img[1880]), .O(
        n14674) );
  MOAI1S U17629 ( .A1(n15780), .A2(n31690), .B1(n13885), .B2(img[856]), .O(
        n14673) );
  NR2 U17630 ( .I1(n14674), .I2(n14673), .O(n14675) );
  ND3 U17631 ( .I1(n14677), .I2(n14676), .I3(n14675), .O(n17158) );
  MOAI1 U17632 ( .A1(n17164), .A2(n13945), .B1(n17158), .B2(n20406), .O(n14702) );
  MOAI1S U17633 ( .A1(n19648), .A2(n31703), .B1(n19642), .B2(img[168]), .O(
        n14678) );
  NR2 U17634 ( .I1(n14679), .I2(n14678), .O(n14682) );
  AOI22S U17635 ( .A1(n15561), .A2(img[1192]), .B1(n13853), .B2(img[1320]), 
        .O(n14681) );
  AOI22S U17636 ( .A1(n18819), .A2(img[40]), .B1(n15657), .B2(img[552]), .O(
        n14680) );
  ND3S U17637 ( .I1(n14682), .I2(n14681), .I3(n14680), .O(n14689) );
  AOI22S U17638 ( .A1(n13865), .A2(img[1832]), .B1(n15630), .B2(img[1576]), 
        .O(n14687) );
  MOAI1S U17639 ( .A1(n13850), .A2(n31624), .B1(n15080), .B2(img[1960]), .O(
        n14684) );
  MOAI1S U17640 ( .A1(n15765), .A2(n31612), .B1(n13837), .B2(img[680]), .O(
        n14683) );
  NR2 U17641 ( .I1(n14684), .I2(n14683), .O(n14686) );
  AOI22S U17642 ( .A1(n19376), .A2(img[808]), .B1(n13845), .B2(img[1448]), .O(
        n14685) );
  ND3S U17643 ( .I1(n14687), .I2(n14686), .I3(n14685), .O(n14688) );
  AOI22S U17644 ( .A1(n13892), .A2(img[1000]), .B1(n15660), .B2(img[232]), .O(
        n14693) );
  AOI22S U17645 ( .A1(n15691), .A2(img[488]), .B1(n15537), .B2(img[360]), .O(
        n14692) );
  AOI22S U17646 ( .A1(n15561), .A2(img[1256]), .B1(n13853), .B2(img[1384]), 
        .O(n14691) );
  AOI22S U17647 ( .A1(n13841), .A2(img[104]), .B1(n13876), .B2(img[616]), .O(
        n14690) );
  AN4S U17648 ( .I1(n14693), .I2(n14692), .I3(n14691), .I4(n14690), .O(n14700)
         );
  MOAI1S U17649 ( .A1(n13850), .A2(n31627), .B1(n15080), .B2(img[2024]), .O(
        n14695) );
  MOAI1S U17650 ( .A1(n15765), .A2(n31615), .B1(n13797), .B2(img[744]), .O(
        n14694) );
  NR2 U17651 ( .I1(n14695), .I2(n14694), .O(n14699) );
  MOAI1S U17652 ( .A1(n15698), .A2(n31623), .B1(n15809), .B2(img[1896]), .O(
        n14697) );
  MOAI1S U17653 ( .A1(n15780), .A2(n31596), .B1(n13886), .B2(img[872]), .O(
        n14696) );
  NR2 U17654 ( .I1(n14697), .I2(n14696), .O(n14698) );
  MOAI1 U17655 ( .A1(n17159), .A2(n16468), .B1(n14706), .B2(n13839), .O(n14701) );
  ND3HT U17656 ( .I1(n14705), .I2(n14704), .I3(n14703), .O(n19573) );
  INV2 U17657 ( .I(n19573), .O(n22942) );
  INV1S U17658 ( .I(n14706), .O(n17161) );
  NR2 U17659 ( .I1(n15448), .I2(n17161), .O(n14708) );
  MOAI1 U17660 ( .A1(n17172), .A2(n17656), .B1(n17173), .B2(n18040), .O(n14707) );
  INV1S U17661 ( .I(n14709), .O(n17179) );
  AOI22S U17662 ( .A1(n13839), .A2(n17166), .B1(n17179), .B2(n13830), .O(
        n14711) );
  AOI22S U17663 ( .A1(n17160), .A2(n13843), .B1(n17178), .B2(n13793), .O(
        n14710) );
  ND3 U17664 ( .I1(n14712), .I2(n14711), .I3(n14710), .O(n14721) );
  MOAI1 U17665 ( .A1(n17164), .A2(n13946), .B1(n17167), .B2(n20439), .O(n14714) );
  MOAI1 U17666 ( .A1(n17159), .A2(n17397), .B1(n17158), .B2(n17938), .O(n14713) );
  NR2 U17667 ( .I1(n14714), .I2(n14713), .O(n14719) );
  AOI22S U17668 ( .A1(n13804), .A2(n17180), .B1(n14715), .B2(n17875), .O(
        n14718) );
  INV1S U17669 ( .I(n14716), .O(n17177) );
  MAOI1S U17670 ( .A1(n17177), .A2(n13846), .B1(n15142), .B2(n17165), .O(
        n14717) );
  ND3 U17671 ( .I1(n14719), .I2(n14718), .I3(n14717), .O(n14720) );
  NR2 U17672 ( .I1(n14721), .I2(n14720), .O(n19575) );
  OR2 U17673 ( .I1(n20969), .I2(n19575), .O(n18484) );
  NR2 U17674 ( .I1(n21728), .I2(n21799), .O(n15371) );
  MOAI1S U17675 ( .A1(n19648), .A2(n31402), .B1(n19642), .B2(img[139]), .O(
        n14722) );
  NR2 U17676 ( .I1(n14723), .I2(n14722), .O(n14726) );
  AOI22S U17677 ( .A1(n13792), .A2(img[1163]), .B1(n15315), .B2(img[1291]), 
        .O(n14725) );
  AOI22S U17678 ( .A1(n13833), .A2(img[11]), .B1(n13876), .B2(img[523]), .O(
        n14724) );
  ND3 U17679 ( .I1(n14726), .I2(n14725), .I3(n14724), .O(n14733) );
  AOI22S U17680 ( .A1(n19036), .A2(img[1803]), .B1(n13874), .B2(img[1547]), 
        .O(n14731) );
  MOAI1S U17681 ( .A1(n13850), .A2(n31418), .B1(n17514), .B2(img[1931]), .O(
        n14728) );
  INV1S U17682 ( .I(n15652), .O(n15343) );
  MOAI1S U17683 ( .A1(n15343), .A2(n31291), .B1(n13797), .B2(img[651]), .O(
        n14727) );
  NR2 U17684 ( .I1(n14728), .I2(n14727), .O(n14730) );
  AOI22S U17685 ( .A1(n19641), .A2(img[779]), .B1(n13845), .B2(img[1419]), .O(
        n14729) );
  ND3S U17686 ( .I1(n14731), .I2(n14730), .I3(n14729), .O(n14732) );
  MOAI1S U17687 ( .A1(n15698), .A2(n31298), .B1(n15080), .B2(img[1995]), .O(
        n14738) );
  INV1S U17688 ( .I(img[1867]), .O(n27355) );
  MOAI1S U17689 ( .A1(n18109), .A2(n27355), .B1(n13885), .B2(img[843]), .O(
        n14737) );
  INV1S U17690 ( .I(img[1739]), .O(n27378) );
  AOI22S U17691 ( .A1(n15799), .A2(img[459]), .B1(n13876), .B2(img[587]), .O(
        n14735) );
  ND2S U17692 ( .I1(n13797), .I2(img[715]), .O(n14734) );
  OAI112HS U17693 ( .C1(n15765), .C2(n27378), .A1(n14735), .B1(n14734), .O(
        n14736) );
  NR3 U17694 ( .I1(n14738), .I2(n14737), .I3(n14736), .O(n14746) );
  INV1S U17695 ( .I(img[1483]), .O(n27688) );
  MOAI1S U17696 ( .A1(n19648), .A2(n31422), .B1(n19642), .B2(img[203]), .O(
        n14740) );
  NR2 U17697 ( .I1(n14741), .I2(n14740), .O(n14745) );
  MOAI1S U17698 ( .A1(n13838), .A2(n31394), .B1(n19290), .B2(img[75]), .O(
        n14743) );
  MOAI1S U17699 ( .A1(n13850), .A2(n31416), .B1(n15315), .B2(img[1355]), .O(
        n14742) );
  NR2 U17700 ( .I1(n14743), .I2(n14742), .O(n14744) );
  ND3 U17701 ( .I1(n14746), .I2(n14745), .I3(n14744), .O(n17665) );
  MOAI1 U17702 ( .A1(n17657), .A2(n13945), .B1(n17665), .B2(n20439), .O(n14821) );
  MOAI1S U17703 ( .A1(n19648), .A2(n31421), .B1(n19642), .B2(img[179]), .O(
        n14747) );
  AOI22S U17704 ( .A1(n15800), .A2(img[1203]), .B1(n15315), .B2(img[1331]), 
        .O(n14750) );
  AOI22S U17705 ( .A1(n19411), .A2(img[51]), .B1(n13876), .B2(img[563]), .O(
        n14749) );
  AOI22S U17706 ( .A1(n13865), .A2(img[1843]), .B1(n20109), .B2(img[1587]), 
        .O(n14756) );
  MOAI1S U17707 ( .A1(n15343), .A2(n31290), .B1(n13898), .B2(img[691]), .O(
        n14752) );
  NR2 U17708 ( .I1(n14753), .I2(n14752), .O(n14755) );
  AOI22S U17709 ( .A1(n13784), .A2(img[819]), .B1(n17862), .B2(img[1459]), .O(
        n14754) );
  ND3 U17710 ( .I1(n14756), .I2(n14755), .I3(n14754), .O(n14757) );
  MOAI1S U17711 ( .A1(n13850), .A2(n31440), .B1(n13896), .B2(img[475]), .O(
        n14764) );
  MOAI1S U17712 ( .A1(n15674), .A2(n31443), .B1(n13876), .B2(img[603]), .O(
        n14763) );
  ND2S U17713 ( .I1(n15800), .I2(img[1243]), .O(n14760) );
  ND2S U17714 ( .I1(n15315), .I2(img[1371]), .O(n14759) );
  ND3S U17715 ( .I1(n14761), .I2(n14760), .I3(n14759), .O(n14762) );
  NR3 U17716 ( .I1(n14764), .I2(n14763), .I3(n14762), .O(n14771) );
  MOAI1S U17717 ( .A1(n15343), .A2(n31367), .B1(n13797), .B2(img[731]), .O(
        n14766) );
  MOAI1S U17718 ( .A1(n15631), .A2(n31463), .B1(n13885), .B2(img[859]), .O(
        n14765) );
  NR2 U17719 ( .I1(n14766), .I2(n14765), .O(n14770) );
  INV1S U17720 ( .I(img[1627]), .O(n27588) );
  MOAI1S U17721 ( .A1(n15698), .A2(n27588), .B1(n20033), .B2(img[2011]), .O(
        n14768) );
  NR2 U17722 ( .I1(n14768), .I2(n14767), .O(n14769) );
  ND3S U17723 ( .I1(n14771), .I2(n14770), .I3(n14769), .O(n17663) );
  MOAI1 U17724 ( .A1(n17659), .A2(n15142), .B1(n17663), .B2(n17931), .O(n14820) );
  MOAI1S U17725 ( .A1(n19648), .A2(n31321), .B1(n19642), .B2(img[171]), .O(
        n14772) );
  NR2 U17726 ( .I1(n14773), .I2(n14772), .O(n14776) );
  AOI22S U17727 ( .A1(n15800), .A2(img[1195]), .B1(n15315), .B2(img[1323]), 
        .O(n14775) );
  AOI22S U17728 ( .A1(n17793), .A2(img[43]), .B1(n13876), .B2(img[555]), .O(
        n14774) );
  ND3 U17729 ( .I1(n14776), .I2(n14775), .I3(n14774), .O(n14783) );
  AOI22S U17730 ( .A1(n13865), .A2(img[1835]), .B1(n15630), .B2(img[1579]), 
        .O(n14781) );
  MOAI1S U17731 ( .A1(n13850), .A2(n31305), .B1(n20193), .B2(img[1963]), .O(
        n14778) );
  MOAI1S U17732 ( .A1(n14914), .A2(n31293), .B1(n13797), .B2(img[683]), .O(
        n14777) );
  NR2 U17733 ( .I1(n14778), .I2(n14777), .O(n14780) );
  ND3S U17734 ( .I1(n14781), .I2(n14780), .I3(n14779), .O(n14782) );
  AOI22S U17735 ( .A1(n15653), .A2(img[931]), .B1(n15773), .B2(img[163]), .O(
        n14787) );
  AOI22S U17736 ( .A1(n15799), .A2(img[419]), .B1(n13800), .B2(img[291]), .O(
        n14786) );
  AOI22S U17737 ( .A1(n15800), .A2(img[1187]), .B1(n15315), .B2(img[1315]), 
        .O(n14785) );
  AOI22S U17738 ( .A1(n18797), .A2(img[35]), .B1(n13876), .B2(img[547]), .O(
        n14784) );
  AN4S U17739 ( .I1(n14787), .I2(n14786), .I3(n14785), .I4(n14784), .O(n14794)
         );
  MOAI1S U17740 ( .A1(n13850), .A2(n31439), .B1(n15080), .B2(img[1955]), .O(
        n14789) );
  MOAI1S U17741 ( .A1(n15343), .A2(n31366), .B1(n13837), .B2(img[675]), .O(
        n14788) );
  NR2 U17742 ( .I1(n14789), .I2(n14788), .O(n14793) );
  MOAI1S U17743 ( .A1(n15698), .A2(n31374), .B1(n15809), .B2(img[1827]), .O(
        n14791) );
  MOAI1S U17744 ( .A1(n15668), .A2(n31458), .B1(n13885), .B2(img[803]), .O(
        n14790) );
  NR2 U17745 ( .I1(n14791), .I2(n14790), .O(n14792) );
  AOI22S U17746 ( .A1(n13880), .A2(img[915]), .B1(n19642), .B2(img[147]), .O(
        n14798) );
  AOI22S U17747 ( .A1(n13859), .A2(img[403]), .B1(n18772), .B2(img[275]), .O(
        n14797) );
  AOI22S U17748 ( .A1(n18922), .A2(img[1171]), .B1(n15315), .B2(img[1299]), 
        .O(n14796) );
  AOI22S U17749 ( .A1(n17515), .A2(img[19]), .B1(n13876), .B2(img[531]), .O(
        n14795) );
  AN4 U17750 ( .I1(n14798), .I2(n14797), .I3(n14796), .I4(n14795), .O(n14805)
         );
  MOAI1S U17751 ( .A1(n13850), .A2(n31308), .B1(n20033), .B2(img[1939]), .O(
        n14800) );
  MOAI1S U17752 ( .A1(n14914), .A2(n31296), .B1(n13898), .B2(img[659]), .O(
        n14799) );
  NR2 U17753 ( .I1(n14800), .I2(n14799), .O(n14804) );
  MOAI1S U17754 ( .A1(n15698), .A2(n31304), .B1(n15809), .B2(img[1811]), .O(
        n14802) );
  MOAI1S U17755 ( .A1(n15668), .A2(n31280), .B1(n13884), .B2(img[787]), .O(
        n14801) );
  NR2 U17756 ( .I1(n14802), .I2(n14801), .O(n14803) );
  ND3P U17757 ( .I1(n14805), .I2(n14804), .I3(n14803), .O(n17662) );
  AOI22S U17758 ( .A1(n17654), .A2(n20124), .B1(n17762), .B2(n17662), .O(
        n14818) );
  AOI22S U17759 ( .A1(n13893), .A2(img[963]), .B1(n15773), .B2(img[195]), .O(
        n14809) );
  AOI22S U17760 ( .A1(n19709), .A2(img[451]), .B1(n18904), .B2(img[323]), .O(
        n14808) );
  AOI22S U17761 ( .A1(n18922), .A2(img[1219]), .B1(n15315), .B2(img[1347]), 
        .O(n14807) );
  AOI22S U17762 ( .A1(n13833), .A2(img[67]), .B1(n13876), .B2(img[579]), .O(
        n14806) );
  INV1S U17763 ( .I(img[1091]), .O(n27615) );
  MOAI1S U17764 ( .A1(n13850), .A2(n27615), .B1(n17617), .B2(img[1987]), .O(
        n14811) );
  MOAI1S U17765 ( .A1(n14914), .A2(n31373), .B1(n13837), .B2(img[707]), .O(
        n14810) );
  NR2 U17766 ( .I1(n14811), .I2(n14810), .O(n14815) );
  MOAI1S U17767 ( .A1(n15698), .A2(n31380), .B1(n15809), .B2(img[1859]), .O(
        n14813) );
  MOAI1S U17768 ( .A1(n15668), .A2(n31355), .B1(n13885), .B2(img[835]), .O(
        n14812) );
  NR2 U17769 ( .I1(n14813), .I2(n14812), .O(n14814) );
  ND3 U17770 ( .I1(n14816), .I2(n14815), .I3(n14814), .O(n17664) );
  ND2S U17771 ( .I1(n17664), .I2(n18040), .O(n14817) );
  OAI112HS U17772 ( .C1(n17655), .C2(n16468), .A1(n14818), .B1(n14817), .O(
        n14819) );
  NR3H U17773 ( .I1(n14821), .I2(n14820), .I3(n14819), .O(n14926) );
  MOAI1S U17774 ( .A1(n13850), .A2(n31381), .B1(n15809), .B2(img[1795]), .O(
        n14824) );
  MOAI1S U17775 ( .A1(n14914), .A2(n31370), .B1(n13837), .B2(img[643]), .O(
        n14823) );
  NR2 U17776 ( .I1(n14824), .I2(n14823), .O(n14827) );
  AOI22S U17777 ( .A1(n19326), .A2(img[771]), .B1(n18751), .B2(img[1411]), .O(
        n14826) );
  AOI22S U17778 ( .A1(n13855), .A2(img[387]), .B1(n15773), .B2(img[131]), .O(
        n14825) );
  ND3S U17779 ( .I1(n14827), .I2(n14826), .I3(n14825), .O(n14834) );
  MOAI1S U17780 ( .A1(n15698), .A2(n31377), .B1(n15786), .B2(img[259]), .O(
        n14829) );
  MOAI1S U17781 ( .A1(n18141), .A2(n31385), .B1(n15657), .B2(img[515]), .O(
        n14828) );
  NR2 U17782 ( .I1(n14829), .I2(n14828), .O(n14832) );
  AOI22S U17783 ( .A1(n13893), .A2(img[899]), .B1(n15315), .B2(img[1283]), .O(
        n14831) );
  AOI22S U17784 ( .A1(n13803), .A2(img[3]), .B1(n15800), .B2(img[1155]), .O(
        n14830) );
  ND3S U17785 ( .I1(n14832), .I2(n14831), .I3(n14830), .O(n14833) );
  NR2 U17786 ( .I1(n14834), .I2(n14833), .O(n17678) );
  AOI22S U17787 ( .A1(n13880), .A2(img[1011]), .B1(n15773), .B2(img[243]), .O(
        n14838) );
  AOI22S U17788 ( .A1(n13879), .A2(img[499]), .B1(n18880), .B2(img[371]), .O(
        n14837) );
  AOI22S U17789 ( .A1(n15800), .A2(img[1267]), .B1(n15315), .B2(img[1395]), 
        .O(n14836) );
  AOI22S U17790 ( .A1(n13803), .A2(img[115]), .B1(n13876), .B2(img[627]), .O(
        n14835) );
  MOAI1S U17791 ( .A1(n13850), .A2(n31417), .B1(n17514), .B2(img[2035]), .O(
        n14840) );
  MOAI1S U17792 ( .A1(n14914), .A2(n31292), .B1(n13797), .B2(img[755]), .O(
        n14839) );
  NR2 U17793 ( .I1(n14840), .I2(n14839), .O(n14844) );
  MOAI1S U17794 ( .A1(n15698), .A2(n31300), .B1(n15809), .B2(img[1907]), .O(
        n14842) );
  MOAI1S U17795 ( .A1(n15780), .A2(n31410), .B1(n15568), .B2(img[883]), .O(
        n14841) );
  NR2 U17796 ( .I1(n14842), .I2(n14841), .O(n14843) );
  ND3 U17797 ( .I1(n14845), .I2(n14844), .I3(n14843), .O(n17680) );
  MOAI1S U17798 ( .A1(n19648), .A2(n31485), .B1(n19642), .B2(img[155]), .O(
        n14846) );
  NR2 U17799 ( .I1(n14847), .I2(n14846), .O(n14850) );
  AOI22S U17800 ( .A1(n15800), .A2(img[1179]), .B1(n15315), .B2(img[1307]), 
        .O(n14849) );
  AOI22S U17801 ( .A1(n13803), .A2(img[27]), .B1(n13876), .B2(img[539]), .O(
        n14848) );
  ND3 U17802 ( .I1(n14850), .I2(n14849), .I3(n14848), .O(n14857) );
  AOI22S U17803 ( .A1(n13863), .A2(img[1819]), .B1(n13874), .B2(img[1563]), 
        .O(n14855) );
  MOAI1S U17804 ( .A1(n13850), .A2(n31437), .B1(n15080), .B2(img[1947]), .O(
        n14852) );
  MOAI1S U17805 ( .A1(n14914), .A2(n31368), .B1(n13898), .B2(img[667]), .O(
        n14851) );
  NR2 U17806 ( .I1(n14852), .I2(n14851), .O(n14854) );
  AOI22S U17807 ( .A1(n19641), .A2(img[795]), .B1(n13845), .B2(img[1435]), .O(
        n14853) );
  ND3 U17808 ( .I1(n14855), .I2(n14854), .I3(n14853), .O(n14856) );
  AOI22S U17809 ( .A1(n13893), .A2(img[995]), .B1(n15773), .B2(img[227]), .O(
        n14861) );
  AOI22S U17810 ( .A1(n13896), .A2(img[483]), .B1(n18995), .B2(img[355]), .O(
        n14860) );
  AOI22S U17811 ( .A1(n15800), .A2(img[1251]), .B1(n13853), .B2(img[1379]), 
        .O(n14859) );
  AOI22S U17812 ( .A1(n20104), .A2(img[99]), .B1(n13876), .B2(img[611]), .O(
        n14858) );
  MOAI1S U17813 ( .A1(n13850), .A2(n31438), .B1(n15080), .B2(img[2019]), .O(
        n14863) );
  MOAI1S U17814 ( .A1(n14914), .A2(n31369), .B1(n13837), .B2(img[739]), .O(
        n14862) );
  NR2 U17815 ( .I1(n14863), .I2(n14862), .O(n14867) );
  MOAI1S U17816 ( .A1(n15698), .A2(n31376), .B1(n15809), .B2(img[1891]), .O(
        n14865) );
  MOAI1S U17817 ( .A1(n15780), .A2(n31457), .B1(n15568), .B2(img[867]), .O(
        n14864) );
  NR2 U17818 ( .I1(n14865), .I2(n14864), .O(n14866) );
  ND3 U17819 ( .I1(n14868), .I2(n14867), .I3(n14866), .O(n17677) );
  MOAI1S U17820 ( .A1(n17675), .A2(n13766), .B1(n17677), .B2(n14869), .O(
        n14870) );
  NR2 U17821 ( .I1(n14871), .I2(n14870), .O(n14925) );
  INV1S U17822 ( .I(img[1147]), .O(n27609) );
  MOAI1S U17823 ( .A1(n13850), .A2(n27609), .B1(n15809), .B2(img[1915]), .O(
        n14873) );
  NR2 U17824 ( .I1(n14873), .I2(n14872), .O(n14876) );
  AOI22S U17825 ( .A1(n15537), .A2(img[379]), .B1(n15773), .B2(img[251]), .O(
        n14874) );
  MOAI1S U17826 ( .A1(n15698), .A2(n31378), .B1(n17514), .B2(img[2043]), .O(
        n14878) );
  MOAI1S U17827 ( .A1(n13789), .A2(n31341), .B1(n13896), .B2(img[507]), .O(
        n14877) );
  NR2 U17828 ( .I1(n14878), .I2(n14877), .O(n14881) );
  AOI22S U17829 ( .A1(n13890), .A2(img[1019]), .B1(n15800), .B2(img[1275]), 
        .O(n14880) );
  AOI22S U17830 ( .A1(n17886), .A2(img[123]), .B1(n13876), .B2(img[635]), .O(
        n14879) );
  ND3S U17831 ( .I1(n14881), .I2(n14880), .I3(n14879), .O(n14882) );
  NR2 U17832 ( .I1(n14883), .I2(n14882), .O(n17670) );
  MOAI1S U17833 ( .A1(n15698), .A2(n31302), .B1(n20033), .B2(img[2003]), .O(
        n14888) );
  MOAI1S U17834 ( .A1(n18109), .A2(n31288), .B1(n15568), .B2(img[851]), .O(
        n14887) );
  AOI22S U17835 ( .A1(n15691), .A2(img[467]), .B1(n13876), .B2(img[595]), .O(
        n14885) );
  ND2S U17836 ( .I1(n13797), .I2(img[723]), .O(n14884) );
  OAI112HS U17837 ( .C1(n15765), .C2(n31294), .A1(n14885), .B1(n14884), .O(
        n14886) );
  NR3 U17838 ( .I1(n14888), .I2(n14887), .I3(n14886), .O(n14895) );
  INV1S U17839 ( .I(img[1491]), .O(n27336) );
  MOAI1S U17840 ( .A1(n15668), .A2(n27336), .B1(n15786), .B2(img[339]), .O(
        n14890) );
  MOAI1S U17841 ( .A1(n13789), .A2(n31267), .B1(n19642), .B2(img[211]), .O(
        n14889) );
  NR2 U17842 ( .I1(n14890), .I2(n14889), .O(n14894) );
  MOAI1S U17843 ( .A1(n13850), .A2(n31306), .B1(n13892), .B2(img[979]), .O(
        n14892) );
  MOAI1S U17844 ( .A1(n13838), .A2(n31263), .B1(n18996), .B2(img[83]), .O(
        n14891) );
  NR2 U17845 ( .I1(n14892), .I2(n14891), .O(n14893) );
  ND3 U17846 ( .I1(n14895), .I2(n14894), .I3(n14893), .O(n17669) );
  MOAI1S U17847 ( .A1(n17670), .A2(n13844), .B1(n17669), .B2(n17938), .O(
        n14923) );
  MOAI1S U17848 ( .A1(n19648), .A2(n31344), .B1(n19642), .B2(img[187]), .O(
        n14897) );
  AOI22S U17849 ( .A1(n13787), .A2(img[1211]), .B1(n13853), .B2(img[1339]), 
        .O(n14900) );
  AOI22S U17850 ( .A1(n13803), .A2(img[59]), .B1(n13876), .B2(img[571]), .O(
        n14899) );
  ND3 U17851 ( .I1(n14901), .I2(n14900), .I3(n14899), .O(n14908) );
  AOI22S U17852 ( .A1(n19215), .A2(img[1851]), .B1(n18837), .B2(img[1595]), 
        .O(n14906) );
  MOAI1S U17853 ( .A1(n13850), .A2(n31382), .B1(n20033), .B2(img[1979]), .O(
        n14903) );
  MOAI1S U17854 ( .A1(n14914), .A2(n31372), .B1(n13797), .B2(img[699]), .O(
        n14902) );
  NR2 U17855 ( .I1(n14903), .I2(n14902), .O(n14905) );
  AOI22S U17856 ( .A1(n13875), .A2(img[827]), .B1(n17827), .B2(img[1467]), .O(
        n14904) );
  ND3S U17857 ( .I1(n14906), .I2(n14905), .I3(n14904), .O(n14907) );
  AOI22S U17858 ( .A1(n15653), .A2(img[1003]), .B1(n15773), .B2(img[235]), .O(
        n14913) );
  AOI22S U17859 ( .A1(n13859), .A2(img[491]), .B1(n18957), .B2(img[363]), .O(
        n14912) );
  AOI22S U17860 ( .A1(n15800), .A2(img[1259]), .B1(n13853), .B2(img[1387]), 
        .O(n14911) );
  AOI22S U17861 ( .A1(n13833), .A2(img[107]), .B1(n13876), .B2(img[619]), .O(
        n14910) );
  MOAI1S U17862 ( .A1(n13850), .A2(n31307), .B1(n15080), .B2(img[2027]), .O(
        n14916) );
  MOAI1S U17863 ( .A1(n14914), .A2(n31295), .B1(n13797), .B2(img[747]), .O(
        n14915) );
  NR2 U17864 ( .I1(n14916), .I2(n14915), .O(n14920) );
  MOAI1S U17865 ( .A1(n15698), .A2(n31303), .B1(n15751), .B2(img[1899]), .O(
        n14918) );
  MOAI1S U17866 ( .A1(n15780), .A2(n31279), .B1(n15568), .B2(img[875]), .O(
        n14917) );
  NR2 U17867 ( .I1(n14918), .I2(n14917), .O(n14919) );
  MOAI1 U17868 ( .A1(n17672), .A2(n17658), .B1(n17671), .B2(n13839), .O(n14922) );
  NR2 U17869 ( .I1(n14923), .I2(n14922), .O(n14924) );
  ND3P U17870 ( .I1(n14926), .I2(n14925), .I3(n14924), .O(n17454) );
  INV2 U17871 ( .I(n13766), .O(n20438) );
  AOI22S U17872 ( .A1(n17664), .A2(n13843), .B1(n20438), .B2(n17654), .O(
        n14928) );
  ND2S U17873 ( .I1(n17665), .I2(n20150), .O(n14927) );
  OAI112HS U17874 ( .C1(n17655), .C2(n17397), .A1(n14928), .B1(n14927), .O(
        n14929) );
  INV1S U17875 ( .I(n17662), .O(n14932) );
  NR2 U17876 ( .I1(n13945), .I2(n14932), .O(n14934) );
  NR2 U17877 ( .I1(n14934), .I2(n14933), .O(n14938) );
  NR2 U17878 ( .I1(n14936), .I2(n14935), .O(n14937) );
  INV1S U17879 ( .I(n19514), .O(n14940) );
  NR2 U17880 ( .I1(n15868), .I2(n21336), .O(n15837) );
  INV1S U17881 ( .I(template_store[44]), .O(n15885) );
  NR2 U17882 ( .I1(n15885), .I2(n15886), .O(n15377) );
  INV1S U17883 ( .I(template_store[42]), .O(n15878) );
  NR2 U17884 ( .I1(n15878), .I2(n15867), .O(n15374) );
  NR2 U17885 ( .I1(n15885), .I2(n21799), .O(n15373) );
  NR2 U17886 ( .I1(n15878), .I2(n21336), .O(n15375) );
  INV1S U17887 ( .I(template_store[40]), .O(n21800) );
  MOAI1S U17888 ( .A1(n19648), .A2(n30925), .B1(n19642), .B2(img[173]), .O(
        n14941) );
  AOI22S U17889 ( .A1(n15561), .A2(img[1197]), .B1(n13853), .B2(img[1325]), 
        .O(n14944) );
  AOI22S U17890 ( .A1(n19411), .A2(img[45]), .B1(n19343), .B2(img[557]), .O(
        n14943) );
  AOI22S U17891 ( .A1(n13865), .A2(img[1837]), .B1(n15630), .B2(img[1581]), 
        .O(n14950) );
  MOAI1S U17892 ( .A1(n13850), .A2(n30883), .B1(n15080), .B2(img[1965]), .O(
        n14947) );
  MOAI1S U17893 ( .A1(n15765), .A2(n30871), .B1(n13797), .B2(img[685]), .O(
        n14946) );
  NR2 U17894 ( .I1(n14947), .I2(n14946), .O(n14949) );
  AOI22S U17895 ( .A1(n13884), .A2(img[813]), .B1(n13845), .B2(img[1453]), .O(
        n14948) );
  ND3S U17896 ( .I1(n14950), .I2(n14949), .I3(n14948), .O(n14951) );
  AOI22S U17897 ( .A1(n15691), .A2(img[509]), .B1(n15800), .B2(img[1277]), .O(
        n14955) );
  ND2S U17898 ( .I1(n17088), .I2(img[1405]), .O(n14954) );
  ND2S U17899 ( .I1(n15657), .I2(img[637]), .O(n14953) );
  ND3S U17900 ( .I1(n14955), .I2(n14954), .I3(n14953), .O(n14959) );
  AOI22S U17901 ( .A1(n15537), .A2(img[381]), .B1(n13803), .B2(img[125]), .O(
        n14957) );
  ND2S U17902 ( .I1(n19642), .I2(img[253]), .O(n14956) );
  OAI112HS U17903 ( .C1(n15698), .C2(n30816), .A1(n14957), .B1(n14956), .O(
        n14958) );
  NR2 U17904 ( .I1(n14959), .I2(n14958), .O(n14966) );
  MOAI1S U17905 ( .A1(n13850), .A2(n30914), .B1(n15080), .B2(img[2045]), .O(
        n14961) );
  MOAI1S U17906 ( .A1(n15765), .A2(n30809), .B1(n13797), .B2(img[765]), .O(
        n14960) );
  NR2 U17907 ( .I1(n14961), .I2(n14960), .O(n14965) );
  MOAI1S U17908 ( .A1(n19648), .A2(n30991), .B1(n13885), .B2(img[893]), .O(
        n14962) );
  NR2 U17909 ( .I1(n14963), .I2(n14962), .O(n14964) );
  MOAI1 U17910 ( .A1(n16706), .A2(n16468), .B1(n16705), .B2(n20969), .O(n15039) );
  MOAI1S U17911 ( .A1(n18141), .A2(n30829), .B1(n15315), .B2(img[1373]), .O(
        n14967) );
  NR2 U17912 ( .I1(n14968), .I2(n14967), .O(n14971) );
  AOI22S U17913 ( .A1(n13893), .A2(img[989]), .B1(n15800), .B2(img[1245]), .O(
        n14970) );
  AOI22S U17914 ( .A1(n18773), .A2(img[93]), .B1(n13876), .B2(img[605]), .O(
        n14969) );
  ND3 U17915 ( .I1(n14971), .I2(n14970), .I3(n14969), .O(n14978) );
  MOAI1S U17916 ( .A1(n15765), .A2(n30811), .B1(n13797), .B2(img[733]), .O(
        n14973) );
  MOAI1S U17917 ( .A1(n15698), .A2(n30818), .B1(n13885), .B2(img[861]), .O(
        n14972) );
  NR2 U17918 ( .I1(n14973), .I2(n14972), .O(n14976) );
  AOI22S U17919 ( .A1(n15537), .A2(img[349]), .B1(n15660), .B2(img[221]), .O(
        n14974) );
  ND3S U17920 ( .I1(n14976), .I2(n14975), .I3(n14974), .O(n14977) );
  AOI22S U17921 ( .A1(n13893), .A2(img[1005]), .B1(n15660), .B2(img[237]), .O(
        n14982) );
  AOI22S U17922 ( .A1(n13859), .A2(img[493]), .B1(n15537), .B2(img[365]), .O(
        n14981) );
  AOI22S U17923 ( .A1(n15561), .A2(img[1261]), .B1(n13853), .B2(img[1389]), 
        .O(n14980) );
  AOI22S U17924 ( .A1(n17335), .A2(img[109]), .B1(n15506), .B2(img[621]), .O(
        n14979) );
  MOAI1S U17925 ( .A1(n13850), .A2(n30885), .B1(n15080), .B2(img[2029]), .O(
        n14984) );
  MOAI1S U17926 ( .A1(n15765), .A2(n30873), .B1(n13797), .B2(img[749]), .O(
        n14983) );
  NR2 U17927 ( .I1(n14984), .I2(n14983), .O(n14988) );
  MOAI1S U17928 ( .A1(n15698), .A2(n30881), .B1(n15809), .B2(img[1901]), .O(
        n14986) );
  MOAI1S U17929 ( .A1(n15668), .A2(n30854), .B1(n13885), .B2(img[877]), .O(
        n14985) );
  NR2 U17930 ( .I1(n14986), .I2(n14985), .O(n14987) );
  ND3 U17931 ( .I1(n14989), .I2(n14988), .I3(n14987), .O(n16707) );
  MOAI1 U17932 ( .A1(n16708), .A2(n20587), .B1(n16707), .B2(n13839), .O(n15038) );
  MOAI1S U17933 ( .A1(n19648), .A2(n30955), .B1(n19642), .B2(img[181]), .O(
        n14990) );
  NR2 U17934 ( .I1(n14991), .I2(n14990), .O(n14994) );
  AOI22S U17935 ( .A1(n15561), .A2(img[1205]), .B1(n13853), .B2(img[1333]), 
        .O(n14993) );
  AOI22S U17936 ( .A1(n18797), .A2(img[53]), .B1(n19343), .B2(img[565]), .O(
        n14992) );
  ND3 U17937 ( .I1(n14994), .I2(n14993), .I3(n14992), .O(n15001) );
  AOI22S U17938 ( .A1(n15809), .A2(img[1845]), .B1(n15630), .B2(img[1589]), 
        .O(n14999) );
  MOAI1S U17939 ( .A1(n13850), .A2(n30941), .B1(n15080), .B2(img[1973]), .O(
        n14996) );
  MOAI1S U17940 ( .A1(n15765), .A2(n30867), .B1(n13837), .B2(img[693]), .O(
        n14995) );
  NR2 U17941 ( .I1(n14996), .I2(n14995), .O(n14998) );
  AOI22S U17942 ( .A1(n13885), .A2(img[821]), .B1(n13845), .B2(img[1461]), .O(
        n14997) );
  ND3S U17943 ( .I1(n14999), .I2(n14998), .I3(n14997), .O(n15000) );
  AOI22S U17944 ( .A1(n15653), .A2(img[901]), .B1(n15660), .B2(img[133]), .O(
        n15005) );
  AOI22S U17945 ( .A1(n13896), .A2(img[389]), .B1(n15537), .B2(img[261]), .O(
        n15004) );
  AOI22S U17946 ( .A1(n15561), .A2(img[1157]), .B1(n13852), .B2(img[1285]), 
        .O(n15003) );
  AOI22S U17947 ( .A1(n17515), .A2(img[5]), .B1(n13876), .B2(img[517]), .O(
        n15002) );
  MOAI1S U17948 ( .A1(n13850), .A2(n30913), .B1(n15080), .B2(img[1925]), .O(
        n15007) );
  MOAI1S U17949 ( .A1(n15765), .A2(n30808), .B1(n13797), .B2(img[645]), .O(
        n15006) );
  NR2 U17950 ( .I1(n15007), .I2(n15006), .O(n15011) );
  MOAI1S U17951 ( .A1(n15698), .A2(n30815), .B1(n13869), .B2(img[1797]), .O(
        n15009) );
  MOAI1S U17952 ( .A1(n15668), .A2(n30908), .B1(n13885), .B2(img[773]), .O(
        n15008) );
  NR2 U17953 ( .I1(n15009), .I2(n15008), .O(n15010) );
  AOI22S U17954 ( .A1(n13892), .A2(img[957]), .B1(n15660), .B2(img[189]), .O(
        n15016) );
  AOI22S U17955 ( .A1(n13859), .A2(img[445]), .B1(n15537), .B2(img[317]), .O(
        n15015) );
  AOI22S U17956 ( .A1(n15561), .A2(img[1213]), .B1(n13853), .B2(img[1341]), 
        .O(n15014) );
  AOI22S U17957 ( .A1(n13833), .A2(img[61]), .B1(n13876), .B2(img[573]), .O(
        n15013) );
  AN4 U17958 ( .I1(n15016), .I2(n15015), .I3(n15014), .I4(n15013), .O(n15023)
         );
  MOAI1S U17959 ( .A1(n13850), .A2(n30915), .B1(n15080), .B2(img[1981]), .O(
        n15018) );
  MOAI1S U17960 ( .A1(n15765), .A2(n30806), .B1(n13837), .B2(img[701]), .O(
        n15017) );
  NR2 U17961 ( .I1(n15018), .I2(n15017), .O(n15022) );
  MOAI1S U17962 ( .A1(n15668), .A2(n30910), .B1(n13885), .B2(img[829]), .O(
        n15019) );
  NR2 U17963 ( .I1(n15020), .I2(n15019), .O(n15021) );
  ND3P U17964 ( .I1(n15023), .I2(n15022), .I3(n15021), .O(n16711) );
  AOI22S U17965 ( .A1(n16712), .A2(n13847), .B1(n17928), .B2(n16711), .O(
        n15036) );
  AOI22S U17966 ( .A1(n16048), .A2(img[909]), .B1(n15660), .B2(img[141]), .O(
        n15027) );
  AOI22S U17967 ( .A1(n13896), .A2(img[397]), .B1(n15537), .B2(img[269]), .O(
        n15026) );
  AOI22S U17968 ( .A1(n15561), .A2(img[1165]), .B1(n13853), .B2(img[1293]), 
        .O(n15025) );
  AOI22S U17969 ( .A1(n17816), .A2(img[13]), .B1(n15506), .B2(img[525]), .O(
        n15024) );
  MOAI1S U17970 ( .A1(n13850), .A2(n30939), .B1(n15080), .B2(img[1933]), .O(
        n15029) );
  MOAI1S U17971 ( .A1(n15765), .A2(n30869), .B1(n13898), .B2(img[653]), .O(
        n15028) );
  NR2 U17972 ( .I1(n15029), .I2(n15028), .O(n15033) );
  MOAI1S U17973 ( .A1(n15698), .A2(n30877), .B1(n15809), .B2(img[1805]), .O(
        n15031) );
  MOAI1S U17974 ( .A1(n15668), .A2(n30961), .B1(n13884), .B2(img[781]), .O(
        n15030) );
  NR2 U17975 ( .I1(n15031), .I2(n15030), .O(n15032) );
  ND3 U17976 ( .I1(n15034), .I2(n15033), .I3(n15032), .O(n16715) );
  ND2S U17977 ( .I1(n16715), .I2(n13830), .O(n15035) );
  NR3HP U17978 ( .I1(n15039), .I2(n15038), .I3(n15037), .O(n15141) );
  MOAI1S U17979 ( .A1(n19648), .A2(n30845), .B1(n19642), .B2(img[149]), .O(
        n15040) );
  AOI22S U17980 ( .A1(n15561), .A2(img[1173]), .B1(n18824), .B2(img[1301]), 
        .O(n15043) );
  AOI22S U17981 ( .A1(n13803), .A2(img[21]), .B1(n13785), .B2(img[533]), .O(
        n15042) );
  ND3 U17982 ( .I1(n15044), .I2(n15043), .I3(n15042), .O(n15051) );
  AOI22S U17983 ( .A1(n13786), .A2(img[1813]), .B1(n15630), .B2(img[1557]), 
        .O(n15049) );
  MOAI1S U17984 ( .A1(n13850), .A2(n30886), .B1(n22928), .B2(img[1941]), .O(
        n15046) );
  MOAI1S U17985 ( .A1(n15765), .A2(n30874), .B1(n13797), .B2(img[661]), .O(
        n15045) );
  NR2 U17986 ( .I1(n15046), .I2(n15045), .O(n15048) );
  AOI22S U17987 ( .A1(n16348), .A2(img[789]), .B1(n13845), .B2(img[1429]), .O(
        n15047) );
  ND3S U17988 ( .I1(n15049), .I2(n15048), .I3(n15047), .O(n15050) );
  NR2P U17989 ( .I1(n15051), .I2(n15050), .O(n16720) );
  MOAI1S U17990 ( .A1(n15698), .A2(n30876), .B1(n15080), .B2(img[1997]), .O(
        n15056) );
  MOAI1S U17991 ( .A1(n15765), .A2(n30868), .B1(n13837), .B2(img[717]), .O(
        n15055) );
  AOI22S U17992 ( .A1(n13828), .A2(img[1869]), .B1(n13885), .B2(img[845]), .O(
        n15053) );
  ND2S U17993 ( .I1(n13879), .I2(img[461]), .O(n15052) );
  OAI112HS U17994 ( .C1(n15668), .C2(n30964), .A1(n15053), .B1(n15052), .O(
        n15054) );
  INV1S U17995 ( .I(img[1229]), .O(n26498) );
  MOAI1S U17996 ( .A1(n13838), .A2(n26498), .B1(n17088), .B2(img[1357]), .O(
        n15058) );
  MOAI1S U17997 ( .A1(n19648), .A2(n30956), .B1(n19642), .B2(img[205]), .O(
        n15057) );
  NR2 U17998 ( .I1(n15058), .I2(n15057), .O(n15062) );
  INV1S U17999 ( .I(img[1101]), .O(n26474) );
  MOAI1S U18000 ( .A1(n13850), .A2(n26474), .B1(n15786), .B2(img[333]), .O(
        n15060) );
  MOAI1S U18001 ( .A1(n15674), .A2(n30947), .B1(n13876), .B2(img[589]), .O(
        n15059) );
  NR2 U18002 ( .I1(n15060), .I2(n15059), .O(n15061) );
  ND3 U18003 ( .I1(n15063), .I2(n15062), .I3(n15061), .O(n16719) );
  MOAI1 U18004 ( .A1(n16720), .A2(n17656), .B1(n16719), .B2(n20439), .O(n15089) );
  MOAI1S U18005 ( .A1(n13850), .A2(n30940), .B1(n22928), .B2(img[2037]), .O(
        n15065) );
  MOAI1S U18006 ( .A1(n15765), .A2(n30870), .B1(n13797), .B2(img[757]), .O(
        n15064) );
  NR2 U18007 ( .I1(n15065), .I2(n15064), .O(n15068) );
  AOI22S U18008 ( .A1(n15537), .A2(img[373]), .B1(n13884), .B2(img[885]), .O(
        n15066) );
  ND3S U18009 ( .I1(n15068), .I2(n15067), .I3(n15066), .O(n15075) );
  MOAI1S U18010 ( .A1(n15668), .A2(n30962), .B1(n13892), .B2(img[1013]), .O(
        n15070) );
  MOAI1S U18011 ( .A1(n15378), .A2(n30976), .B1(n13876), .B2(img[629]), .O(
        n15069) );
  NR2 U18012 ( .I1(n15070), .I2(n15069), .O(n15073) );
  AOI22S U18013 ( .A1(n17515), .A2(img[117]), .B1(n15315), .B2(img[1397]), .O(
        n15072) );
  AOI22S U18014 ( .A1(n13855), .A2(img[501]), .B1(n15800), .B2(img[1269]), .O(
        n15071) );
  ND3 U18015 ( .I1(n15073), .I2(n15072), .I3(n15071), .O(n15074) );
  NR2P U18016 ( .I1(n15075), .I2(n15074), .O(n16722) );
  AOI22S U18017 ( .A1(n13893), .A2(img[981]), .B1(n15660), .B2(img[213]), .O(
        n15079) );
  AOI22S U18018 ( .A1(n13896), .A2(img[469]), .B1(n15537), .B2(img[341]), .O(
        n15078) );
  AOI22S U18019 ( .A1(n15561), .A2(img[1237]), .B1(n17088), .B2(img[1365]), 
        .O(n15077) );
  AOI22S U18020 ( .A1(n18983), .A2(img[85]), .B1(n13876), .B2(img[597]), .O(
        n15076) );
  MOAI1S U18021 ( .A1(n13850), .A2(n30884), .B1(n15080), .B2(img[2005]), .O(
        n15082) );
  MOAI1S U18022 ( .A1(n15765), .A2(n30872), .B1(n13898), .B2(img[725]), .O(
        n15081) );
  NR2 U18023 ( .I1(n15082), .I2(n15081), .O(n15086) );
  MOAI1S U18024 ( .A1(n15698), .A2(n30880), .B1(n15809), .B2(img[1877]), .O(
        n15084) );
  MOAI1S U18025 ( .A1(n15780), .A2(n30853), .B1(n15568), .B2(img[853]), .O(
        n15083) );
  NR2 U18026 ( .I1(n15084), .I2(n15083), .O(n15085) );
  ND3 U18027 ( .I1(n15087), .I2(n15086), .I3(n15085), .O(n16721) );
  MOAI1 U18028 ( .A1(n16722), .A2(n13947), .B1(n16721), .B2(n17938), .O(n15088) );
  MOAI1S U18029 ( .A1(n19648), .A2(n30786), .B1(n19642), .B2(img[157]), .O(
        n15090) );
  AOI22S U18030 ( .A1(n15561), .A2(img[1181]), .B1(n18963), .B2(img[1309]), 
        .O(n15093) );
  AOI22S U18031 ( .A1(n20104), .A2(img[29]), .B1(n13876), .B2(img[541]), .O(
        n15092) );
  INV1S U18032 ( .I(n16758), .O(n16064) );
  AOI22S U18033 ( .A1(n13863), .A2(img[1821]), .B1(n15630), .B2(img[1565]), 
        .O(n15099) );
  MOAI1S U18034 ( .A1(n13850), .A2(n30822), .B1(n22928), .B2(img[1949]), .O(
        n15096) );
  MOAI1S U18035 ( .A1(n15765), .A2(n30812), .B1(n13898), .B2(img[669]), .O(
        n15095) );
  NR2 U18036 ( .I1(n15096), .I2(n15095), .O(n15098) );
  AOI22S U18037 ( .A1(n17835), .A2(img[797]), .B1(n13845), .B2(img[1437]), .O(
        n15097) );
  ND3S U18038 ( .I1(n15099), .I2(n15098), .I3(n15097), .O(n15100) );
  NR2P U18039 ( .I1(n15101), .I2(n15100), .O(n16725) );
  AOI22S U18040 ( .A1(n13893), .A2(img[965]), .B1(n17088), .B2(img[1349]), .O(
        n15105) );
  AOI22S U18041 ( .A1(n13896), .A2(img[453]), .B1(n15537), .B2(img[325]), .O(
        n15104) );
  AOI22S U18042 ( .A1(n17335), .A2(img[69]), .B1(n15800), .B2(img[1221]), .O(
        n15103) );
  AOI22S U18043 ( .A1(n19215), .A2(img[1861]), .B1(n15660), .B2(img[197]), .O(
        n15102) );
  AN4S U18044 ( .I1(n15105), .I2(n15104), .I3(n15103), .I4(n15102), .O(n15112)
         );
  MOAI1S U18045 ( .A1(n15765), .A2(n30807), .B1(n13837), .B2(img[709]), .O(
        n15107) );
  MOAI1S U18046 ( .A1(n13850), .A2(n30916), .B1(n13876), .B2(img[581]), .O(
        n15106) );
  NR2 U18047 ( .I1(n15107), .I2(n15106), .O(n15111) );
  INV1S U18048 ( .I(img[1605]), .O(n26150) );
  MOAI1S U18049 ( .A1(n15698), .A2(n26150), .B1(n22928), .B2(img[1989]), .O(
        n15109) );
  MOAI1S U18050 ( .A1(n15780), .A2(n30911), .B1(n13884), .B2(img[837]), .O(
        n15108) );
  NR2 U18051 ( .I1(n15109), .I2(n15108), .O(n15110) );
  MOAI1 U18052 ( .A1(n16725), .A2(n13766), .B1(n16727), .B2(n18040), .O(n15138) );
  MOAI1S U18053 ( .A1(n19648), .A2(n30999), .B1(n19642), .B2(img[165]), .O(
        n15114) );
  NR2 U18054 ( .I1(n15115), .I2(n15114), .O(n15118) );
  AOI22S U18055 ( .A1(n15561), .A2(img[1189]), .B1(n18910), .B2(img[1317]), 
        .O(n15117) );
  AOI22S U18056 ( .A1(n19290), .A2(img[37]), .B1(n13825), .B2(img[549]), .O(
        n15116) );
  ND3 U18057 ( .I1(n15118), .I2(n15117), .I3(n15116), .O(n15125) );
  AOI22S U18058 ( .A1(n19023), .A2(img[1829]), .B1(n15630), .B2(img[1573]), 
        .O(n15123) );
  MOAI1S U18059 ( .A1(n13850), .A2(n30820), .B1(n22928), .B2(img[1957]), .O(
        n15120) );
  AOI22S U18060 ( .A1(n13885), .A2(img[805]), .B1(n13845), .B2(img[1445]), .O(
        n15121) );
  ND3S U18061 ( .I1(n15123), .I2(n15122), .I3(n15121), .O(n15124) );
  NR2P U18062 ( .I1(n15125), .I2(n15124), .O(n16728) );
  AOI22S U18063 ( .A1(n13893), .A2(img[997]), .B1(n15660), .B2(img[229]), .O(
        n15129) );
  AOI22S U18064 ( .A1(n15799), .A2(img[485]), .B1(n15537), .B2(img[357]), .O(
        n15128) );
  AOI22S U18065 ( .A1(n15561), .A2(img[1253]), .B1(n17088), .B2(img[1381]), 
        .O(n15127) );
  AOI22S U18066 ( .A1(n18797), .A2(img[101]), .B1(n13883), .B2(img[613]), .O(
        n15126) );
  MOAI1S U18067 ( .A1(n13850), .A2(n30823), .B1(n22928), .B2(img[2021]), .O(
        n15131) );
  MOAI1S U18068 ( .A1(n15765), .A2(n30813), .B1(n13898), .B2(img[741]), .O(
        n15130) );
  NR2 U18069 ( .I1(n15131), .I2(n15130), .O(n15135) );
  INV1S U18070 ( .I(img[1637]), .O(n26166) );
  MOAI1S U18071 ( .A1(n15698), .A2(n26166), .B1(n15809), .B2(img[1893]), .O(
        n15133) );
  INV1S U18072 ( .I(img[1509]), .O(n26092) );
  MOAI1S U18073 ( .A1(n15668), .A2(n26092), .B1(n15568), .B2(img[869]), .O(
        n15132) );
  NR2 U18074 ( .I1(n15133), .I2(n15132), .O(n15134) );
  MOAI1 U18075 ( .A1(n16728), .A2(n17397), .B1(n16729), .B2(n21062), .O(n15137) );
  NR2P U18076 ( .I1(n15138), .I2(n15137), .O(n15139) );
  ND3HT U18077 ( .I1(n15141), .I2(n15140), .I3(n15139), .O(n21245) );
  OAI22S U18078 ( .A1(n16713), .A2(n16468), .B1(n16722), .B2(n19462), .O(
        n15146) );
  ND2S U18079 ( .I1(n16729), .I2(n17931), .O(n15144) );
  ND2S U18080 ( .I1(n16715), .I2(n13847), .O(n15143) );
  OAI112HS U18081 ( .C1(n16706), .C2(n17397), .A1(n15144), .B1(n15143), .O(
        n15145) );
  INV1S U18082 ( .I(n16719), .O(n15148) );
  MOAI1 U18083 ( .A1(n15148), .A2(n20421), .B1(n16705), .B2(n13846), .O(n15151) );
  INV1S U18084 ( .I(n16707), .O(n15149) );
  MOAI1 U18085 ( .A1(n15149), .A2(n15448), .B1(n16727), .B2(n13843), .O(n15150) );
  NR2 U18086 ( .I1(n15151), .I2(n15150), .O(n15155) );
  INV1S U18087 ( .I(n19495), .O(n15157) );
  NR2 U18088 ( .I1(n21800), .I2(n21726), .O(n15600) );
  INV1S U18089 ( .I(template_store[41]), .O(n15875) );
  OAI22S U18090 ( .A1(n31979), .A2(n19648), .B1(n15378), .B2(n31981), .O(
        n15159) );
  NR2 U18091 ( .I1(n15159), .I2(n15158), .O(n15162) );
  AOI22S U18092 ( .A1(n15800), .A2(img[1276]), .B1(n17088), .B2(img[1404]), 
        .O(n15161) );
  AOI22S U18093 ( .A1(n17864), .A2(img[124]), .B1(n13876), .B2(img[636]), .O(
        n15160) );
  ND3 U18094 ( .I1(n15162), .I2(n15161), .I3(n15160), .O(n15169) );
  MOAI1S U18095 ( .A1(n13850), .A2(n31856), .B1(n15080), .B2(img[2044]), .O(
        n15164) );
  MOAI1S U18096 ( .A1(n15806), .A2(n31844), .B1(n13797), .B2(img[764]), .O(
        n15163) );
  NR2 U18097 ( .I1(n15164), .I2(n15163), .O(n15167) );
  AOI22S U18098 ( .A1(n13865), .A2(img[1916]), .B1(n18837), .B2(img[1660]), 
        .O(n15166) );
  AOI22S U18099 ( .A1(n13884), .A2(img[892]), .B1(n13845), .B2(img[1532]), .O(
        n15165) );
  NR2 U18100 ( .I1(n15169), .I2(n15168), .O(n17916) );
  AOI22S U18101 ( .A1(n13893), .A2(img[900]), .B1(n19642), .B2(img[132]), .O(
        n15173) );
  AOI22S U18102 ( .A1(n15799), .A2(img[388]), .B1(n15786), .B2(img[260]), .O(
        n15172) );
  AOI22S U18103 ( .A1(n15800), .A2(img[1156]), .B1(n13824), .B2(img[1284]), 
        .O(n15171) );
  AOI22S U18104 ( .A1(n13841), .A2(img[4]), .B1(n13876), .B2(img[516]), .O(
        n15170) );
  MOAI1S U18105 ( .A1(n13850), .A2(n31855), .B1(n20193), .B2(img[1924]), .O(
        n15175) );
  MOAI1S U18106 ( .A1(n15806), .A2(n31843), .B1(n13797), .B2(img[644]), .O(
        n15174) );
  NR2 U18107 ( .I1(n15175), .I2(n15174), .O(n15179) );
  MOAI1S U18108 ( .A1(n15698), .A2(n31851), .B1(n15809), .B2(img[1796]), .O(
        n15177) );
  MOAI1S U18109 ( .A1(n15780), .A2(n31825), .B1(n13885), .B2(img[772]), .O(
        n15176) );
  NR2 U18110 ( .I1(n15177), .I2(n15176), .O(n15178) );
  ND3 U18111 ( .I1(n15180), .I2(n15179), .I3(n15178), .O(n17915) );
  OAI22S U18112 ( .A1(n31902), .A2(n19648), .B1(n15378), .B2(n31904), .O(
        n15182) );
  NR2 U18113 ( .I1(n15182), .I2(n15181), .O(n15185) );
  AOI22S U18114 ( .A1(n15800), .A2(img[1196]), .B1(n13824), .B2(img[1324]), 
        .O(n15184) );
  AOI22S U18115 ( .A1(n20104), .A2(img[44]), .B1(n15657), .B2(img[556]), .O(
        n15183) );
  ND3S U18116 ( .I1(n15185), .I2(n15184), .I3(n15183), .O(n15192) );
  MOAI1S U18117 ( .A1(n13850), .A2(n31894), .B1(n20033), .B2(img[1964]), .O(
        n15187) );
  MOAI1S U18118 ( .A1(n15806), .A2(n31777), .B1(n13797), .B2(img[684]), .O(
        n15186) );
  NR2 U18119 ( .I1(n15187), .I2(n15186), .O(n15190) );
  AOI22S U18120 ( .A1(n13863), .A2(img[1836]), .B1(n18837), .B2(img[1580]), 
        .O(n15189) );
  AOI22S U18121 ( .A1(n15568), .A2(img[812]), .B1(n13845), .B2(img[1452]), .O(
        n15188) );
  ND3S U18122 ( .I1(n15190), .I2(n15189), .I3(n15188), .O(n15191) );
  NR2 U18123 ( .I1(n15192), .I2(n15191), .O(n17918) );
  AOI22S U18124 ( .A1(n13893), .A2(img[908]), .B1(n19642), .B2(img[140]), .O(
        n15196) );
  AOI22S U18125 ( .A1(n15799), .A2(img[396]), .B1(n15786), .B2(img[268]), .O(
        n15195) );
  AOI22S U18126 ( .A1(n15800), .A2(img[1164]), .B1(n17088), .B2(img[1292]), 
        .O(n15194) );
  AOI22S U18127 ( .A1(n17793), .A2(img[12]), .B1(n18681), .B2(img[524]), .O(
        n15193) );
  AN4S U18128 ( .I1(n15196), .I2(n15195), .I3(n15194), .I4(n15193), .O(n15203)
         );
  MOAI1S U18129 ( .A1(n13850), .A2(n31793), .B1(n15080), .B2(img[1932]), .O(
        n15198) );
  MOAI1S U18130 ( .A1(n15806), .A2(n31781), .B1(n13837), .B2(img[652]), .O(
        n15197) );
  NR2 U18131 ( .I1(n15198), .I2(n15197), .O(n15202) );
  MOAI1S U18132 ( .A1(n15698), .A2(n31789), .B1(n15809), .B2(img[1804]), .O(
        n15200) );
  MOAI1S U18133 ( .A1(n15780), .A2(n31762), .B1(n15568), .B2(img[780]), .O(
        n15199) );
  ND3 U18134 ( .I1(n15203), .I2(n15202), .I3(n15201), .O(n17917) );
  MOAI1 U18135 ( .A1(n17918), .A2(n16468), .B1(n17917), .B2(n13830), .O(n15252) );
  MOAI1S U18136 ( .A1(n13850), .A2(n31857), .B1(n17382), .B2(img[1604]), .O(
        n15205) );
  MOAI1S U18137 ( .A1(n15806), .A2(n31845), .B1(n13898), .B2(img[708]), .O(
        n15204) );
  NR2 U18138 ( .I1(n15205), .I2(n15204), .O(n15208) );
  AOI22S U18139 ( .A1(n13882), .A2(img[452]), .B1(n15751), .B2(img[1860]), .O(
        n15207) );
  AOI22S U18140 ( .A1(n15660), .A2(img[196]), .B1(n15568), .B2(img[836]), .O(
        n15206) );
  ND3S U18141 ( .I1(n15208), .I2(n15207), .I3(n15206), .O(n15215) );
  MOAI1S U18142 ( .A1(n13838), .A2(n31811), .B1(n14909), .B2(img[68]), .O(
        n15209) );
  NR2 U18143 ( .I1(n15210), .I2(n15209), .O(n15213) );
  AOI22S U18144 ( .A1(n15537), .A2(img[324]), .B1(n13827), .B2(img[1348]), .O(
        n15212) );
  AOI22S U18145 ( .A1(n13893), .A2(img[964]), .B1(n15506), .B2(img[580]), .O(
        n15211) );
  ND3S U18146 ( .I1(n15213), .I2(n15212), .I3(n15211), .O(n15214) );
  NR2 U18147 ( .I1(n15215), .I2(n15214), .O(n17924) );
  AOI22S U18148 ( .A1(n19403), .A2(img[932]), .B1(n19642), .B2(img[164]), .O(
        n15219) );
  AOI22S U18149 ( .A1(n13882), .A2(img[420]), .B1(n18831), .B2(img[292]), .O(
        n15218) );
  AOI22S U18150 ( .A1(n15800), .A2(img[1188]), .B1(n17088), .B2(img[1316]), 
        .O(n15217) );
  AOI22S U18151 ( .A1(n13833), .A2(img[36]), .B1(n13825), .B2(img[548]), .O(
        n15216) );
  AN4 U18152 ( .I1(n15219), .I2(n15218), .I3(n15217), .I4(n15216), .O(n15226)
         );
  MOAI1S U18153 ( .A1(n13850), .A2(n31915), .B1(n22928), .B2(img[1956]), .O(
        n15221) );
  MOAI1S U18154 ( .A1(n15806), .A2(n31839), .B1(n13898), .B2(img[676]), .O(
        n15220) );
  NR2 U18155 ( .I1(n15221), .I2(n15220), .O(n15225) );
  MOAI1S U18156 ( .A1(n15780), .A2(n31933), .B1(n13884), .B2(img[804]), .O(
        n15222) );
  NR2 U18157 ( .I1(n15223), .I2(n15222), .O(n15224) );
  ND3P U18158 ( .I1(n15226), .I2(n15225), .I3(n15224), .O(n17920) );
  AOI22S U18159 ( .A1(n15653), .A2(img[924]), .B1(n15773), .B2(img[156]), .O(
        n15230) );
  AOI22S U18160 ( .A1(n13882), .A2(img[412]), .B1(n19710), .B2(img[284]), .O(
        n15229) );
  AOI22S U18161 ( .A1(n15652), .A2(img[1692]), .B1(n13837), .B2(img[668]), .O(
        n15228) );
  AOI22S U18162 ( .A1(n15630), .A2(img[1564]), .B1(n13788), .B2(img[1052]), 
        .O(n15227) );
  MOAI1S U18163 ( .A1(n13872), .A2(n31943), .B1(n13801), .B2(img[28]), .O(
        n15232) );
  MOAI1S U18164 ( .A1(n13790), .A2(n31931), .B1(n15800), .B2(img[1180]), .O(
        n15231) );
  NR2 U18165 ( .I1(n15232), .I2(n15231), .O(n15236) );
  MOAI1S U18166 ( .A1(n15668), .A2(n31935), .B1(n15080), .B2(img[1948]), .O(
        n15234) );
  MOAI1S U18167 ( .A1(n15277), .A2(n31927), .B1(n15809), .B2(img[1820]), .O(
        n15233) );
  NR2 U18168 ( .I1(n15234), .I2(n15233), .O(n15235) );
  ND3 U18169 ( .I1(n15237), .I2(n15236), .I3(n15235), .O(n17919) );
  AOI22S U18170 ( .A1(n17920), .A2(n20124), .B1(n20438), .B2(n17919), .O(
        n15250) );
  AOI22S U18171 ( .A1(n16048), .A2(img[1012]), .B1(n15315), .B2(img[1396]), 
        .O(n15241) );
  AOI22S U18172 ( .A1(n22928), .A2(img[2036]), .B1(n13825), .B2(img[628]), .O(
        n15240) );
  AOI22S U18173 ( .A1(n15537), .A2(img[372]), .B1(n19642), .B2(img[244]), .O(
        n15239) );
  AOI22S U18174 ( .A1(n18819), .A2(img[116]), .B1(n15800), .B2(img[1268]), .O(
        n15238) );
  AN4S U18175 ( .I1(n15241), .I2(n15240), .I3(n15239), .I4(n15238), .O(n15248)
         );
  MOAI1S U18176 ( .A1(n15698), .A2(n31790), .B1(n15809), .B2(img[1908]), .O(
        n15243) );
  MOAI1S U18177 ( .A1(n15806), .A2(n31782), .B1(n13797), .B2(img[756]), .O(
        n15242) );
  NR2 U18178 ( .I1(n15243), .I2(n15242), .O(n15247) );
  MOAI1S U18179 ( .A1(n15668), .A2(n31763), .B1(n13879), .B2(img[500]), .O(
        n15245) );
  MOAI1S U18180 ( .A1(n13850), .A2(n31794), .B1(n15568), .B2(img[884]), .O(
        n15244) );
  NR2 U18181 ( .I1(n15245), .I2(n15244), .O(n15246) );
  ND3 U18182 ( .I1(n15248), .I2(n15247), .I3(n15246), .O(n17921) );
  ND2S U18183 ( .I1(n17921), .I2(n13846), .O(n15249) );
  OAI112HS U18184 ( .C1(n17924), .C2(n20421), .A1(n15250), .B1(n15249), .O(
        n15251) );
  NR3H U18185 ( .I1(n15253), .I2(n15252), .I3(n15251), .O(n15355) );
  MOAI1S U18186 ( .A1(n18141), .A2(n31799), .B1(n13879), .B2(img[404]), .O(
        n15255) );
  MOAI1S U18187 ( .A1(n13838), .A2(n31873), .B1(n19024), .B2(img[1556]), .O(
        n15254) );
  NR2 U18188 ( .I1(n15255), .I2(n15254), .O(n15258) );
  AOI22S U18189 ( .A1(n13890), .A2(img[916]), .B1(n13783), .B2(img[1300]), .O(
        n15257) );
  AOI22S U18190 ( .A1(n18983), .A2(img[20]), .B1(n13876), .B2(img[532]), .O(
        n15256) );
  ND3 U18191 ( .I1(n15258), .I2(n15257), .I3(n15256), .O(n15265) );
  MOAI1S U18192 ( .A1(n15343), .A2(n31779), .B1(n13898), .B2(img[660]), .O(
        n15259) );
  NR2 U18193 ( .I1(n15260), .I2(n15259), .O(n15263) );
  AOI22S U18194 ( .A1(n13884), .A2(img[788]), .B1(n17862), .B2(img[1428]), .O(
        n15262) );
  AOI22S U18195 ( .A1(n15537), .A2(img[276]), .B1(n19642), .B2(img[148]), .O(
        n15261) );
  ND3S U18196 ( .I1(n15263), .I2(n15262), .I3(n15261), .O(n15264) );
  AOI22S U18197 ( .A1(n13893), .A2(img[948]), .B1(n15773), .B2(img[180]), .O(
        n15269) );
  AOI22S U18198 ( .A1(n13882), .A2(img[436]), .B1(n18995), .B2(img[308]), .O(
        n15268) );
  AOI22S U18199 ( .A1(n15800), .A2(img[1204]), .B1(n17088), .B2(img[1332]), 
        .O(n15267) );
  AOI22S U18200 ( .A1(n18983), .A2(img[52]), .B1(n13876), .B2(img[564]), .O(
        n15266) );
  MOAI1S U18201 ( .A1(n13850), .A2(n31795), .B1(n22928), .B2(img[1972]), .O(
        n15271) );
  MOAI1S U18202 ( .A1(n15343), .A2(n31783), .B1(n13837), .B2(img[692]), .O(
        n15270) );
  NR2 U18203 ( .I1(n15271), .I2(n15270), .O(n15275) );
  MOAI1S U18204 ( .A1(n15698), .A2(n31791), .B1(n15809), .B2(img[1844]), .O(
        n15273) );
  MOAI1S U18205 ( .A1(n15780), .A2(n31764), .B1(n13884), .B2(img[820]), .O(
        n15272) );
  NR2 U18206 ( .I1(n15273), .I2(n15272), .O(n15274) );
  ND3 U18207 ( .I1(n15276), .I2(n15275), .I3(n15274), .O(n17929) );
  MOAI1 U18208 ( .A1(n17930), .A2(n17656), .B1(n17929), .B2(n14174), .O(n15302) );
  MOAI1S U18209 ( .A1(n18109), .A2(n31834), .B1(n22928), .B2(img[2020]), .O(
        n15279) );
  MOAI1S U18210 ( .A1(n15277), .A2(n31928), .B1(n18837), .B2(img[1636]), .O(
        n15278) );
  NR2 U18211 ( .I1(n15279), .I2(n15278), .O(n15282) );
  AOI22S U18212 ( .A1(n13893), .A2(img[996]), .B1(n15800), .B2(img[1252]), .O(
        n15281) );
  AOI22S U18213 ( .A1(n15537), .A2(img[356]), .B1(n18911), .B2(img[1124]), .O(
        n15280) );
  ND3S U18214 ( .I1(n15282), .I2(n15281), .I3(n15280), .O(n15289) );
  MOAI1S U18215 ( .A1(n15378), .A2(n31938), .B1(n13879), .B2(img[484]), .O(
        n15284) );
  NR2 U18216 ( .I1(n15284), .I2(n15283), .O(n15287) );
  AOI22S U18217 ( .A1(n15652), .A2(img[1764]), .B1(n13837), .B2(img[740]), .O(
        n15286) );
  AOI22S U18218 ( .A1(n13841), .A2(img[100]), .B1(n13876), .B2(img[612]), .O(
        n15285) );
  NR2 U18219 ( .I1(n15289), .I2(n15288), .O(n17933) );
  AOI22S U18220 ( .A1(n13860), .A2(img[980]), .B1(n19642), .B2(img[212]), .O(
        n15293) );
  AOI22S U18221 ( .A1(n13882), .A2(img[468]), .B1(n19710), .B2(img[340]), .O(
        n15292) );
  AOI22S U18222 ( .A1(n15800), .A2(img[1236]), .B1(n15315), .B2(img[1364]), 
        .O(n15291) );
  AOI22S U18223 ( .A1(n18797), .A2(img[84]), .B1(n13876), .B2(img[596]), .O(
        n15290) );
  MOAI1S U18224 ( .A1(n13850), .A2(n31895), .B1(n20193), .B2(img[2004]), .O(
        n15295) );
  MOAI1S U18225 ( .A1(n15343), .A2(n31778), .B1(n13837), .B2(img[724]), .O(
        n15294) );
  NR2 U18226 ( .I1(n15295), .I2(n15294), .O(n15299) );
  MOAI1S U18227 ( .A1(n15698), .A2(n31786), .B1(n15809), .B2(img[1876]), .O(
        n15297) );
  MOAI1S U18228 ( .A1(n15780), .A2(n31888), .B1(n13885), .B2(img[852]), .O(
        n15296) );
  NR2 U18229 ( .I1(n15297), .I2(n15296), .O(n15298) );
  ND3 U18230 ( .I1(n15300), .I2(n15299), .I3(n15298), .O(n17932) );
  MOAI1 U18231 ( .A1(n17933), .A2(n15448), .B1(n17932), .B2(n17938), .O(n15301) );
  OAI22S U18232 ( .A1(n31818), .A2(n19648), .B1(n15378), .B2(n31820), .O(
        n15304) );
  NR2 U18233 ( .I1(n15304), .I2(n15303), .O(n15307) );
  AOI22S U18234 ( .A1(n13802), .A2(img[1212]), .B1(n17088), .B2(img[1340]), 
        .O(n15306) );
  AOI22S U18235 ( .A1(n13833), .A2(img[60]), .B1(n13876), .B2(img[572]), .O(
        n15305) );
  ND3S U18236 ( .I1(n15307), .I2(n15306), .I3(n15305), .O(n15314) );
  MOAI1S U18237 ( .A1(n13850), .A2(n31858), .B1(n22928), .B2(img[1980]), .O(
        n15309) );
  MOAI1S U18238 ( .A1(n15343), .A2(n31846), .B1(n13837), .B2(img[700]), .O(
        n15308) );
  NR2 U18239 ( .I1(n15309), .I2(n15308), .O(n15312) );
  AOI22S U18240 ( .A1(n13863), .A2(img[1852]), .B1(n13874), .B2(img[1596]), 
        .O(n15311) );
  AOI22S U18241 ( .A1(n15568), .A2(img[828]), .B1(n13845), .B2(img[1468]), .O(
        n15310) );
  ND3S U18242 ( .I1(n15312), .I2(n15311), .I3(n15310), .O(n15313) );
  NR2 U18243 ( .I1(n15314), .I2(n15313), .O(n17937) );
  AOI22S U18244 ( .A1(n13892), .A2(img[1004]), .B1(n19642), .B2(img[236]), .O(
        n15319) );
  AOI22S U18245 ( .A1(n13882), .A2(img[492]), .B1(n15786), .B2(img[364]), .O(
        n15318) );
  AOI22S U18246 ( .A1(n15800), .A2(img[1260]), .B1(n15315), .B2(img[1388]), 
        .O(n15317) );
  AOI22S U18247 ( .A1(n17778), .A2(img[108]), .B1(n13876), .B2(img[620]), .O(
        n15316) );
  MOAI1S U18248 ( .A1(n13850), .A2(n31897), .B1(n22928), .B2(img[2028]), .O(
        n15321) );
  MOAI1S U18249 ( .A1(n15343), .A2(n31780), .B1(n13797), .B2(img[748]), .O(
        n15320) );
  NR2 U18250 ( .I1(n15321), .I2(n15320), .O(n15325) );
  INV1S U18251 ( .I(n18297), .O(n20038) );
  MOAI1S U18252 ( .A1(n15780), .A2(n31890), .B1(n13885), .B2(img[876]), .O(
        n15322) );
  MOAI1 U18253 ( .A1(n17937), .A2(n17658), .B1(n17936), .B2(n13839), .O(n15352) );
  OAI22S U18254 ( .A1(n31963), .A2(n19648), .B1(n15378), .B2(n31965), .O(
        n15328) );
  NR2 U18255 ( .I1(n15328), .I2(n15327), .O(n15331) );
  AOI22S U18256 ( .A1(n18909), .A2(img[1244]), .B1(n13824), .B2(img[1372]), 
        .O(n15330) );
  AOI22S U18257 ( .A1(n18797), .A2(img[92]), .B1(n15506), .B2(img[604]), .O(
        n15329) );
  ND3S U18258 ( .I1(n15331), .I2(n15330), .I3(n15329), .O(n15338) );
  MOAI1S U18259 ( .A1(n13850), .A2(n31916), .B1(n15080), .B2(img[2012]), .O(
        n15333) );
  MOAI1S U18260 ( .A1(n15343), .A2(n31840), .B1(n13797), .B2(img[732]), .O(
        n15332) );
  NR2 U18261 ( .I1(n15333), .I2(n15332), .O(n15336) );
  AOI22S U18262 ( .A1(n15809), .A2(img[1884]), .B1(n13874), .B2(img[1628]), 
        .O(n15335) );
  AOI22S U18263 ( .A1(n13884), .A2(img[860]), .B1(n17862), .B2(img[1500]), .O(
        n15334) );
  ND3S U18264 ( .I1(n15336), .I2(n15335), .I3(n15334), .O(n15337) );
  NR2 U18265 ( .I1(n15338), .I2(n15337), .O(n17940) );
  AOI22S U18266 ( .A1(n16048), .A2(img[972]), .B1(n15773), .B2(img[204]), .O(
        n15342) );
  AOI22S U18267 ( .A1(n13896), .A2(img[460]), .B1(n18831), .B2(img[332]), .O(
        n15341) );
  AOI22S U18268 ( .A1(n15800), .A2(img[1228]), .B1(n13854), .B2(img[1356]), 
        .O(n15340) );
  AOI22S U18269 ( .A1(n13801), .A2(img[76]), .B1(n13876), .B2(img[588]), .O(
        n15339) );
  MOAI1S U18270 ( .A1(n13850), .A2(n31796), .B1(n22928), .B2(img[1996]), .O(
        n15345) );
  MOAI1S U18271 ( .A1(n15343), .A2(n31784), .B1(n13898), .B2(img[716]), .O(
        n15344) );
  NR2 U18272 ( .I1(n15345), .I2(n15344), .O(n15349) );
  MOAI1S U18273 ( .A1(n15698), .A2(n31792), .B1(n19215), .B2(img[1868]), .O(
        n15347) );
  MOAI1S U18274 ( .A1(n15780), .A2(n31765), .B1(n13884), .B2(img[844]), .O(
        n15346) );
  NR2 U18275 ( .I1(n15347), .I2(n15346), .O(n15348) );
  ND3 U18276 ( .I1(n15350), .I2(n15349), .I3(n15348), .O(n17939) );
  MOAI1 U18277 ( .A1(n17940), .A2(n20587), .B1(n17939), .B2(n20439), .O(n15351) );
  NR2P U18278 ( .I1(n15352), .I2(n15351), .O(n15353) );
  ND3P U18279 ( .I1(n15355), .I2(n15354), .I3(n15353), .O(n15356) );
  INV1S U18280 ( .I(n17939), .O(n15357) );
  NR2 U18281 ( .I1(n20421), .I2(n15357), .O(n15362) );
  OAI22S U18282 ( .A1(n17916), .A2(n13947), .B1(n17918), .B2(n17397), .O(
        n15361) );
  AOI22S U18283 ( .A1(n17917), .A2(n13847), .B1(n20438), .B2(n17920), .O(
        n15359) );
  ND2S U18284 ( .I1(n17919), .I2(n17762), .O(n15358) );
  OAI112HS U18285 ( .C1(n17924), .C2(n18196), .A1(n15359), .B1(n15358), .O(
        n15360) );
  NR3 U18286 ( .I1(n15362), .I2(n15361), .I3(n15360), .O(n15370) );
  INV1S U18287 ( .I(n17921), .O(n15363) );
  NR2 U18288 ( .I1(n15365), .I2(n15364), .O(n15369) );
  OAI22S U18289 ( .A1(n17933), .A2(n20587), .B1(n17937), .B2(n15142), .O(
        n15366) );
  NR2 U18290 ( .I1(n15367), .I2(n15366), .O(n15368) );
  AOI13HS U18291 ( .B1(n15370), .B2(n15369), .B3(n15368), .A1(n20969), .O(
        n19602) );
  AO12 U18292 ( .B1(n22927), .B2(n20863), .A1(n19602), .O(n20711) );
  INV2 U18293 ( .I(n20711), .O(n21231) );
  NR2 U18294 ( .I1(n15875), .I2(n21231), .O(n15599) );
  HA1 U18295 ( .A(n15372), .B(n15371), .C(n15838), .S(n15598) );
  NR2 U18296 ( .I1(n21800), .I2(n21231), .O(n15850) );
  NR2 U18297 ( .I1(n15868), .I2(n15886), .O(n15849) );
  HA1 U18298 ( .A(n15374), .B(n15373), .C(n15376), .S(n15848) );
  MOAI1S U18299 ( .A1(n13894), .A2(n30523), .B1(n13892), .B2(img[918]), .O(
        n15380) );
  MOAI1S U18300 ( .A1(n15378), .A2(n30519), .B1(n15506), .B2(img[534]), .O(
        n15379) );
  NR2 U18301 ( .I1(n15380), .I2(n15379), .O(n15383) );
  AOI22S U18302 ( .A1(n13803), .A2(img[22]), .B1(n15315), .B2(img[1302]), .O(
        n15382) );
  AOI22S U18303 ( .A1(n13786), .A2(img[1814]), .B1(n15800), .B2(img[1174]), 
        .O(n15381) );
  ND3S U18304 ( .I1(n15383), .I2(n15382), .I3(n15381), .O(n15390) );
  AOI22S U18305 ( .A1(n13845), .A2(img[1430]), .B1(n15630), .B2(img[1558]), 
        .O(n15388) );
  MOAI1S U18306 ( .A1(n13850), .A2(n30490), .B1(n22928), .B2(img[1942]), .O(
        n15385) );
  MOAI1S U18307 ( .A1(n15765), .A2(n30381), .B1(n13837), .B2(img[662]), .O(
        n15384) );
  NR2 U18308 ( .I1(n15385), .I2(n15384), .O(n15387) );
  AOI22S U18309 ( .A1(n15537), .A2(img[278]), .B1(n13885), .B2(img[790]), .O(
        n15386) );
  ND3S U18310 ( .I1(n15388), .I2(n15387), .I3(n15386), .O(n15389) );
  AOI22S U18311 ( .A1(n13892), .A2(img[1006]), .B1(n15660), .B2(img[238]), .O(
        n15394) );
  AOI22S U18312 ( .A1(n13858), .A2(img[494]), .B1(n15537), .B2(img[366]), .O(
        n15393) );
  AOI22S U18313 ( .A1(n15561), .A2(img[1262]), .B1(n15315), .B2(img[1390]), 
        .O(n15392) );
  AOI22S U18314 ( .A1(n17886), .A2(img[110]), .B1(n13785), .B2(img[622]), .O(
        n15391) );
  MOAI1S U18315 ( .A1(n13850), .A2(n30491), .B1(n22928), .B2(img[2030]), .O(
        n15396) );
  MOAI1S U18316 ( .A1(n15765), .A2(n30382), .B1(n13898), .B2(img[750]), .O(
        n15395) );
  NR2 U18317 ( .I1(n15396), .I2(n15395), .O(n15400) );
  MOAI1S U18318 ( .A1(n15698), .A2(n30390), .B1(n13870), .B2(img[1902]), .O(
        n15398) );
  MOAI1S U18319 ( .A1(n15780), .A2(n30487), .B1(n13886), .B2(img[878]), .O(
        n15397) );
  NR2 U18320 ( .I1(n15398), .I2(n15397), .O(n15399) );
  ND3P U18321 ( .I1(n15401), .I2(n15400), .I3(n15399), .O(n16477) );
  MOAI1 U18322 ( .A1(n16471), .A2(n17656), .B1(n16477), .B2(n13839), .O(n15475) );
  MOAI1S U18323 ( .A1(n15698), .A2(n30387), .B1(n15809), .B2(img[1838]), .O(
        n15403) );
  MOAI1S U18324 ( .A1(n15765), .A2(n30379), .B1(n13898), .B2(img[686]), .O(
        n15402) );
  NR2 U18325 ( .I1(n15403), .I2(n15402), .O(n15406) );
  AOI22S U18326 ( .A1(n15691), .A2(img[430]), .B1(n19326), .B2(img[814]), .O(
        n15405) );
  AOI22S U18327 ( .A1(n15537), .A2(img[302]), .B1(n15660), .B2(img[174]), .O(
        n15404) );
  ND3S U18328 ( .I1(n15406), .I2(n15405), .I3(n15404), .O(n15413) );
  AOI22S U18329 ( .A1(n13845), .A2(img[1454]), .B1(n18988), .B2(img[1070]), 
        .O(n15411) );
  MOAI1S U18330 ( .A1(n15674), .A2(n30497), .B1(n13876), .B2(img[558]), .O(
        n15408) );
  MOAI1S U18331 ( .A1(n19648), .A2(n30503), .B1(n15800), .B2(img[1198]), .O(
        n15407) );
  NR2 U18332 ( .I1(n15408), .I2(n15407), .O(n15410) );
  AOI22S U18333 ( .A1(n22928), .A2(img[1966]), .B1(n18963), .B2(img[1326]), 
        .O(n15409) );
  ND3S U18334 ( .I1(n15411), .I2(n15410), .I3(n15409), .O(n15412) );
  AOI22S U18335 ( .A1(n13892), .A2(img[950]), .B1(n15660), .B2(img[182]), .O(
        n15417) );
  AOI22S U18336 ( .A1(n15691), .A2(img[438]), .B1(n15537), .B2(img[310]), .O(
        n15416) );
  AOI22S U18337 ( .A1(n15561), .A2(img[1206]), .B1(n13854), .B2(img[1334]), 
        .O(n15415) );
  AOI22S U18338 ( .A1(n17335), .A2(img[54]), .B1(n20102), .B2(img[566]), .O(
        n15414) );
  MOAI1S U18339 ( .A1(n13850), .A2(n30395), .B1(n22928), .B2(img[1974]), .O(
        n15419) );
  MOAI1S U18340 ( .A1(n15765), .A2(n30383), .B1(n13837), .B2(img[694]), .O(
        n15418) );
  NR2 U18341 ( .I1(n15419), .I2(n15418), .O(n15423) );
  MOAI1S U18342 ( .A1(n15698), .A2(n30391), .B1(n18885), .B2(img[1846]), .O(
        n15421) );
  MOAI1S U18343 ( .A1(n15780), .A2(n30364), .B1(n13886), .B2(img[822]), .O(
        n15420) );
  NR2 U18344 ( .I1(n15421), .I2(n15420), .O(n15422) );
  ND3 U18345 ( .I1(n15424), .I2(n15423), .I3(n15422), .O(n16474) );
  MOAI1 U18346 ( .A1(n16491), .A2(n16468), .B1(n16474), .B2(n14174), .O(n15474) );
  MOAI1S U18347 ( .A1(n19648), .A2(n30475), .B1(n19642), .B2(img[134]), .O(
        n15425) );
  NR2 U18348 ( .I1(n15426), .I2(n15425), .O(n15429) );
  AOI22S U18349 ( .A1(n15561), .A2(img[1158]), .B1(n15315), .B2(img[1286]), 
        .O(n15428) );
  AOI22S U18350 ( .A1(n17515), .A2(img[6]), .B1(n15506), .B2(img[518]), .O(
        n15427) );
  ND3S U18351 ( .I1(n15429), .I2(n15428), .I3(n15427), .O(n15436) );
  AOI22S U18352 ( .A1(n19036), .A2(img[1798]), .B1(n15630), .B2(img[1542]), 
        .O(n15434) );
  MOAI1S U18353 ( .A1(n13850), .A2(n30332), .B1(n22928), .B2(img[1926]), .O(
        n15431) );
  MOAI1S U18354 ( .A1(n15765), .A2(n30320), .B1(n13797), .B2(img[646]), .O(
        n15430) );
  NR2 U18355 ( .I1(n15431), .I2(n15430), .O(n15433) );
  AOI22S U18356 ( .A1(n13885), .A2(img[774]), .B1(n13845), .B2(img[1414]), .O(
        n15432) );
  ND3S U18357 ( .I1(n15434), .I2(n15433), .I3(n15432), .O(n15435) );
  NR2 U18358 ( .I1(n15436), .I2(n15435), .O(n16466) );
  AOI22S U18359 ( .A1(n15653), .A2(img[998]), .B1(n15660), .B2(img[230]), .O(
        n15440) );
  AOI22S U18360 ( .A1(n15691), .A2(img[486]), .B1(n15537), .B2(img[358]), .O(
        n15439) );
  AOI22S U18361 ( .A1(n15561), .A2(img[1254]), .B1(n17088), .B2(img[1382]), 
        .O(n15438) );
  AOI22S U18362 ( .A1(n17335), .A2(img[102]), .B1(n15506), .B2(img[614]), .O(
        n15437) );
  MOAI1S U18363 ( .A1(n13850), .A2(n30436), .B1(n22928), .B2(img[2022]), .O(
        n15442) );
  MOAI1S U18364 ( .A1(n15765), .A2(n30319), .B1(n13837), .B2(img[742]), .O(
        n15441) );
  NR2 U18365 ( .I1(n15442), .I2(n15441), .O(n15446) );
  MOAI1S U18366 ( .A1(n15698), .A2(n30327), .B1(n15809), .B2(img[1894]), .O(
        n15444) );
  MOAI1S U18367 ( .A1(n15668), .A2(n30429), .B1(n13885), .B2(img[870]), .O(
        n15443) );
  NR2 U18368 ( .I1(n15444), .I2(n15443), .O(n15445) );
  ND3 U18369 ( .I1(n15447), .I2(n15446), .I3(n15445), .O(n16470) );
  AOI22S U18370 ( .A1(n16048), .A2(img[982]), .B1(n15660), .B2(img[214]), .O(
        n15452) );
  AOI22S U18371 ( .A1(n13859), .A2(img[470]), .B1(n15537), .B2(img[342]), .O(
        n15451) );
  AOI22S U18372 ( .A1(n15561), .A2(img[1238]), .B1(n17088), .B2(img[1366]), 
        .O(n15450) );
  AOI22S U18373 ( .A1(n13833), .A2(img[86]), .B1(n13785), .B2(img[598]), .O(
        n15449) );
  AN4 U18374 ( .I1(n15452), .I2(n15451), .I3(n15450), .I4(n15449), .O(n15459)
         );
  MOAI1S U18375 ( .A1(n13850), .A2(n30492), .B1(n22928), .B2(img[2006]), .O(
        n15454) );
  MOAI1S U18376 ( .A1(n15765), .A2(n30380), .B1(n13837), .B2(img[726]), .O(
        n15453) );
  NR2 U18377 ( .I1(n15454), .I2(n15453), .O(n15458) );
  MOAI1S U18378 ( .A1(n15668), .A2(n30488), .B1(n15568), .B2(img[854]), .O(
        n15455) );
  NR2 U18379 ( .I1(n15456), .I2(n15455), .O(n15457) );
  ND3 U18380 ( .I1(n15459), .I2(n15458), .I3(n15457), .O(n16475) );
  AOI22S U18381 ( .A1(n16470), .A2(n19483), .B1(n17938), .B2(n16475), .O(
        n15472) );
  AOI22S U18382 ( .A1(n13892), .A2(img[934]), .B1(n15660), .B2(img[166]), .O(
        n15463) );
  AOI22S U18383 ( .A1(n15691), .A2(img[422]), .B1(n15537), .B2(img[294]), .O(
        n15462) );
  AOI22S U18384 ( .A1(n15561), .A2(img[1190]), .B1(n17088), .B2(img[1318]), 
        .O(n15461) );
  AOI22S U18385 ( .A1(n13801), .A2(img[38]), .B1(n13876), .B2(img[550]), .O(
        n15460) );
  MOAI1S U18386 ( .A1(n13850), .A2(n30434), .B1(n22928), .B2(img[1958]), .O(
        n15465) );
  MOAI1S U18387 ( .A1(n15765), .A2(n30316), .B1(n13797), .B2(img[678]), .O(
        n15464) );
  NR2 U18388 ( .I1(n15465), .I2(n15464), .O(n15469) );
  MOAI1S U18389 ( .A1(n15780), .A2(n30427), .B1(n13886), .B2(img[806]), .O(
        n15466) );
  NR2 U18390 ( .I1(n15467), .I2(n15466), .O(n15468) );
  ND2S U18391 ( .I1(n16465), .I2(n20613), .O(n15471) );
  OAI112HS U18392 ( .C1(n16466), .C2(n13946), .A1(n15472), .B1(n15471), .O(
        n15473) );
  MOAI1S U18393 ( .A1(n13850), .A2(n30333), .B1(n22928), .B2(img[2046]), .O(
        n15477) );
  MOAI1S U18394 ( .A1(n15765), .A2(n30321), .B1(n13837), .B2(img[766]), .O(
        n15476) );
  NR2 U18395 ( .I1(n15477), .I2(n15476), .O(n15480) );
  MAOI1S U18396 ( .A1(n19252), .A2(img[894]), .B1(n30329), .B2(n15698), .O(
        n15479) );
  ND3S U18397 ( .I1(n15480), .I2(n15479), .I3(n15478), .O(n15487) );
  MOAI1S U18398 ( .A1(n13838), .A2(n30287), .B1(n13896), .B2(img[510]), .O(
        n15481) );
  NR2 U18399 ( .I1(n15482), .I2(n15481), .O(n15485) );
  AOI22S U18400 ( .A1(n13893), .A2(img[1022]), .B1(n17323), .B2(img[1406]), 
        .O(n15484) );
  AOI22S U18401 ( .A1(n19411), .A2(img[126]), .B1(n13876), .B2(img[638]), .O(
        n15483) );
  NR2P U18402 ( .I1(n15487), .I2(n15486), .O(n16488) );
  AOI22S U18403 ( .A1(n13880), .A2(img[990]), .B1(n15660), .B2(img[222]), .O(
        n15491) );
  AOI22S U18404 ( .A1(n15691), .A2(img[478]), .B1(n15537), .B2(img[350]), .O(
        n15490) );
  AOI22S U18405 ( .A1(n15561), .A2(img[1246]), .B1(n18975), .B2(img[1374]), 
        .O(n15489) );
  AOI22S U18406 ( .A1(n19290), .A2(img[94]), .B1(n15506), .B2(img[606]), .O(
        n15488) );
  MOAI1S U18407 ( .A1(n13850), .A2(n30435), .B1(n22928), .B2(img[2014]), .O(
        n15493) );
  MOAI1S U18408 ( .A1(n15765), .A2(n30317), .B1(n13898), .B2(img[734]), .O(
        n15492) );
  NR2 U18409 ( .I1(n15493), .I2(n15492), .O(n15497) );
  MOAI1S U18410 ( .A1(n15698), .A2(n30325), .B1(n19023), .B2(img[1886]), .O(
        n15495) );
  MOAI1S U18411 ( .A1(n15668), .A2(n30428), .B1(n13886), .B2(img[862]), .O(
        n15494) );
  NR2 U18412 ( .I1(n15495), .I2(n15494), .O(n15496) );
  ND3 U18413 ( .I1(n15498), .I2(n15497), .I3(n15496), .O(n16493) );
  MOAI1 U18414 ( .A1(n16488), .A2(n13844), .B1(n16493), .B2(n20406), .O(n15524) );
  MOAI1S U18415 ( .A1(n15698), .A2(n30393), .B1(n22928), .B2(img[1934]), .O(
        n15500) );
  MOAI1S U18416 ( .A1(n15765), .A2(n30385), .B1(n13797), .B2(img[654]), .O(
        n15499) );
  NR2 U18417 ( .I1(n15500), .I2(n15499), .O(n15503) );
  AOI22S U18418 ( .A1(n15660), .A2(img[142]), .B1(n13845), .B2(img[1422]), .O(
        n15502) );
  AOI22S U18419 ( .A1(n15691), .A2(img[398]), .B1(n15751), .B2(img[1806]), .O(
        n15501) );
  ND3S U18420 ( .I1(n15503), .I2(n15502), .I3(n15501), .O(n15511) );
  MOAI1S U18421 ( .A1(n13850), .A2(n30397), .B1(n15800), .B2(img[1166]), .O(
        n15505) );
  MOAI1S U18422 ( .A1(n15674), .A2(n30346), .B1(n13884), .B2(img[782]), .O(
        n15504) );
  NR2 U18423 ( .I1(n15505), .I2(n15504), .O(n15509) );
  AOI22S U18424 ( .A1(n15537), .A2(img[270]), .B1(n17277), .B2(img[1294]), .O(
        n15508) );
  AOI22S U18425 ( .A1(n13861), .A2(img[910]), .B1(n15506), .B2(img[526]), .O(
        n15507) );
  ND3S U18426 ( .I1(n15509), .I2(n15508), .I3(n15507), .O(n15510) );
  AOI22S U18427 ( .A1(n16048), .A2(img[974]), .B1(n15660), .B2(img[206]), .O(
        n15515) );
  AOI22S U18428 ( .A1(n15691), .A2(img[462]), .B1(n15537), .B2(img[334]), .O(
        n15514) );
  AOI22S U18429 ( .A1(n15561), .A2(img[1230]), .B1(n13853), .B2(img[1358]), 
        .O(n15513) );
  AOI22S U18430 ( .A1(n13803), .A2(img[78]), .B1(n13876), .B2(img[590]), .O(
        n15512) );
  MOAI1S U18431 ( .A1(n13850), .A2(n30396), .B1(n22928), .B2(img[1998]), .O(
        n15517) );
  MOAI1S U18432 ( .A1(n15765), .A2(n30384), .B1(n13797), .B2(img[718]), .O(
        n15516) );
  NR2 U18433 ( .I1(n15517), .I2(n15516), .O(n15521) );
  MOAI1S U18434 ( .A1(n15698), .A2(n30392), .B1(n20038), .B2(img[1870]), .O(
        n15519) );
  MOAI1S U18435 ( .A1(n15668), .A2(n30365), .B1(n15568), .B2(img[846]), .O(
        n15518) );
  NR2 U18436 ( .I1(n15519), .I2(n15518), .O(n15520) );
  MOAI1 U18437 ( .A1(n16482), .A2(n13945), .B1(n16476), .B2(n20263), .O(n15523) );
  NR2 U18438 ( .I1(n15524), .I2(n15523), .O(n15577) );
  MOAI1S U18439 ( .A1(n19648), .A2(n30420), .B1(n19642), .B2(img[158]), .O(
        n15525) );
  AOI22S U18440 ( .A1(n15561), .A2(img[1182]), .B1(n18778), .B2(img[1310]), 
        .O(n15528) );
  AOI22S U18441 ( .A1(n13833), .A2(img[30]), .B1(n13876), .B2(img[542]), .O(
        n15527) );
  ND3 U18442 ( .I1(n15529), .I2(n15528), .I3(n15527), .O(n15536) );
  AOI22S U18443 ( .A1(n19036), .A2(img[1822]), .B1(n15630), .B2(img[1566]), 
        .O(n15534) );
  MOAI1S U18444 ( .A1(n13850), .A2(n30437), .B1(n22928), .B2(img[1950]), .O(
        n15531) );
  MOAI1S U18445 ( .A1(n15765), .A2(n30318), .B1(n13837), .B2(img[670]), .O(
        n15530) );
  NR2 U18446 ( .I1(n15531), .I2(n15530), .O(n15533) );
  AOI22S U18447 ( .A1(n13885), .A2(img[798]), .B1(n13845), .B2(img[1438]), .O(
        n15532) );
  ND3S U18448 ( .I1(n15534), .I2(n15533), .I3(n15532), .O(n15535) );
  NR2P U18449 ( .I1(n15536), .I2(n15535), .O(n16485) );
  AOI22S U18450 ( .A1(n16048), .A2(img[1014]), .B1(n15660), .B2(img[246]), .O(
        n15541) );
  AOI22S U18451 ( .A1(n15799), .A2(img[502]), .B1(n15537), .B2(img[374]), .O(
        n15540) );
  AOI22S U18452 ( .A1(n15561), .A2(img[1270]), .B1(n17088), .B2(img[1398]), 
        .O(n15539) );
  AOI22S U18453 ( .A1(n19411), .A2(img[118]), .B1(n13785), .B2(img[630]), .O(
        n15538) );
  AN4S U18454 ( .I1(n15541), .I2(n15540), .I3(n15539), .I4(n15538), .O(n15548)
         );
  MOAI1S U18455 ( .A1(n13850), .A2(n30398), .B1(n22928), .B2(img[2038]), .O(
        n15543) );
  MOAI1S U18456 ( .A1(n15765), .A2(n30386), .B1(n13837), .B2(img[758]), .O(
        n15542) );
  NR2 U18457 ( .I1(n15543), .I2(n15542), .O(n15547) );
  MOAI1S U18458 ( .A1(n15698), .A2(n30394), .B1(n13870), .B2(img[1910]), .O(
        n15545) );
  MOAI1S U18459 ( .A1(n15668), .A2(n30367), .B1(n13885), .B2(img[886]), .O(
        n15544) );
  NR2 U18460 ( .I1(n15545), .I2(n15544), .O(n15546) );
  MOAI1 U18461 ( .A1(n16485), .A2(n13766), .B1(n16481), .B2(n13846), .O(n15575) );
  MOAI1S U18462 ( .A1(n19648), .A2(n30294), .B1(n15773), .B2(img[190]), .O(
        n15549) );
  AOI22S U18463 ( .A1(n15561), .A2(img[1214]), .B1(n17088), .B2(img[1342]), 
        .O(n15552) );
  AOI22S U18464 ( .A1(n18819), .A2(img[62]), .B1(n19343), .B2(img[574]), .O(
        n15551) );
  ND3 U18465 ( .I1(n15553), .I2(n15552), .I3(n15551), .O(n15560) );
  AOI22S U18466 ( .A1(n19023), .A2(img[1854]), .B1(n20109), .B2(img[1598]), 
        .O(n15558) );
  MOAI1S U18467 ( .A1(n13850), .A2(n30334), .B1(n22928), .B2(img[1982]), .O(
        n15555) );
  MOAI1S U18468 ( .A1(n15765), .A2(n30322), .B1(n13797), .B2(img[702]), .O(
        n15554) );
  NR2 U18469 ( .I1(n15555), .I2(n15554), .O(n15557) );
  AOI22S U18470 ( .A1(n13885), .A2(img[830]), .B1(n13845), .B2(img[1470]), .O(
        n15556) );
  NR2P U18471 ( .I1(n15560), .I2(n15559), .O(n16483) );
  AOI22S U18472 ( .A1(n15653), .A2(img[966]), .B1(n15773), .B2(img[198]), .O(
        n15565) );
  AOI22S U18473 ( .A1(n13896), .A2(img[454]), .B1(n18982), .B2(img[326]), .O(
        n15564) );
  AOI22S U18474 ( .A1(n15561), .A2(img[1222]), .B1(n18789), .B2(img[1350]), 
        .O(n15563) );
  AOI22S U18475 ( .A1(n13801), .A2(img[70]), .B1(n15506), .B2(img[582]), .O(
        n15562) );
  AN4 U18476 ( .I1(n15565), .I2(n15564), .I3(n15563), .I4(n15562), .O(n15573)
         );
  MOAI1S U18477 ( .A1(n13850), .A2(n30335), .B1(n22928), .B2(img[1990]), .O(
        n15567) );
  MOAI1S U18478 ( .A1(n15765), .A2(n30323), .B1(n13797), .B2(img[710]), .O(
        n15566) );
  NR2 U18479 ( .I1(n15567), .I2(n15566), .O(n15572) );
  MOAI1S U18480 ( .A1(n15698), .A2(n30331), .B1(n15751), .B2(img[1862]), .O(
        n15570) );
  MOAI1S U18481 ( .A1(n15780), .A2(n30305), .B1(n15568), .B2(img[838]), .O(
        n15569) );
  NR2 U18482 ( .I1(n15570), .I2(n15569), .O(n15571) );
  ND3 U18483 ( .I1(n15573), .I2(n15572), .I3(n15571), .O(n16490) );
  MOAI1 U18484 ( .A1(n16483), .A2(n17658), .B1(n16490), .B2(n18040), .O(n15574) );
  NR2 U18485 ( .I1(n15575), .I2(n15574), .O(n15576) );
  ND2F U18486 ( .I1(n21254), .I2(n20809), .O(n29513) );
  ND2S U18487 ( .I1(n16490), .I2(n13843), .O(n15582) );
  ND2S U18488 ( .I1(n16470), .I2(n17931), .O(n15581) );
  ND2S U18489 ( .I1(n16475), .I2(n20263), .O(n15580) );
  ND3S U18490 ( .I1(n15582), .I2(n15581), .I3(n15580), .O(n15586) );
  AOI22S U18491 ( .A1(n16465), .A2(n13804), .B1(n21062), .B2(n16477), .O(
        n15584) );
  ND2S U18492 ( .I1(n16474), .I2(n17875), .O(n15583) );
  OAI112HS U18493 ( .C1(n16471), .C2(n13945), .A1(n15584), .B1(n15583), .O(
        n15585) );
  NR2 U18494 ( .I1(n15586), .I2(n15585), .O(n15593) );
  MOAI1S U18495 ( .A1(n16482), .A2(n13946), .B1(n16481), .B2(n13839), .O(
        n15588) );
  OAI22S U18496 ( .A1(n16485), .A2(n17656), .B1(n16483), .B2(n15142), .O(
        n15587) );
  NR2 U18497 ( .I1(n15588), .I2(n15587), .O(n15592) );
  NR2 U18498 ( .I1(n15590), .I2(n15589), .O(n15591) );
  INV1S U18499 ( .I(n19474), .O(n15594) );
  NR2 U18500 ( .I1(n15875), .I2(n21729), .O(n15906) );
  NR2 U18501 ( .I1(n15885), .I2(n21336), .O(n15905) );
  NR2 U18502 ( .I1(n15875), .I2(n21726), .O(n15597) );
  NR2 U18503 ( .I1(n15878), .I2(n21231), .O(n15596) );
  NR2 U18504 ( .I1(n15885), .I2(n15867), .O(n15836) );
  INV1S U18505 ( .I(template_store[46]), .O(n21730) );
  NR2 U18506 ( .I1(n21730), .I2(n21799), .O(n15835) );
  NR2 U18507 ( .I1(n21800), .I2(n21729), .O(n15842) );
  NR2 U18508 ( .I1(n15878), .I2(n21726), .O(n15903) );
  MOAI1S U18509 ( .A1(n15698), .A2(n30146), .B1(n15809), .B2(img[1799]), .O(
        n15602) );
  MOAI1S U18510 ( .A1(n15765), .A2(n30138), .B1(n13898), .B2(img[647]), .O(
        n15601) );
  NR2 U18511 ( .I1(n15602), .I2(n15601), .O(n15605) );
  AOI22S U18512 ( .A1(n16348), .A2(img[775]), .B1(n13845), .B2(img[1415]), .O(
        n15604) );
  AOI22S U18513 ( .A1(n15691), .A2(img[391]), .B1(n15660), .B2(img[135]), .O(
        n15603) );
  ND3S U18514 ( .I1(n15605), .I2(n15604), .I3(n15603), .O(n15612) );
  MOAI1S U18515 ( .A1(n13850), .A2(n30190), .B1(n13841), .B2(img[7]), .O(
        n15607) );
  MOAI1 U18516 ( .A1(n18141), .A2(n30158), .B1(n15786), .B2(img[263]), .O(
        n15606) );
  NR2 U18517 ( .I1(n15607), .I2(n15606), .O(n15610) );
  AOI22S U18518 ( .A1(n15653), .A2(img[903]), .B1(n13824), .B2(img[1287]), .O(
        n15609) );
  AOI22S U18519 ( .A1(n13787), .A2(img[1159]), .B1(n13876), .B2(img[519]), .O(
        n15608) );
  MOAI1S U18520 ( .A1(n15765), .A2(n30141), .B1(n13797), .B2(img[735]), .O(
        n15616) );
  AOI22S U18521 ( .A1(n13882), .A2(img[479]), .B1(n13884), .B2(img[863]), .O(
        n15614) );
  ND2S U18522 ( .I1(n15653), .I2(img[991]), .O(n15613) );
  OAI112HS U18523 ( .C1(n15668), .C2(n30122), .A1(n15614), .B1(n15613), .O(
        n15615) );
  MOAI1S U18524 ( .A1(n13790), .A2(n30110), .B1(n15657), .B2(img[607]), .O(
        n15619) );
  MOAI1S U18525 ( .A1(n13838), .A2(n30106), .B1(n19642), .B2(img[223]), .O(
        n15618) );
  NR2 U18526 ( .I1(n15619), .I2(n15618), .O(n15623) );
  MOAI1S U18527 ( .A1(n13850), .A2(n30153), .B1(n22928), .B2(img[2015]), .O(
        n15621) );
  MOAI1S U18528 ( .A1(n15631), .A2(n30241), .B1(n14909), .B2(img[95]), .O(
        n15620) );
  NR2 U18529 ( .I1(n15621), .I2(n15620), .O(n15622) );
  ND3 U18530 ( .I1(n15624), .I2(n15623), .I3(n15622), .O(n16229) );
  MOAI1 U18531 ( .A1(n16230), .A2(n13946), .B1(n16229), .B2(n17931), .O(n15708) );
  MOAI1S U18532 ( .A1(n13850), .A2(n30091), .B1(n15080), .B2(img[1975]), .O(
        n15626) );
  MOAI1S U18533 ( .A1(n18109), .A2(n30071), .B1(n13885), .B2(img[823]), .O(
        n15625) );
  NR2 U18534 ( .I1(n15626), .I2(n15625), .O(n15629) );
  AOI22S U18535 ( .A1(n13837), .A2(img[695]), .B1(n15652), .B2(img[1719]), .O(
        n15628) );
  AOI22S U18536 ( .A1(n15653), .A2(img[951]), .B1(n17816), .B2(img[55]), .O(
        n15627) );
  ND3S U18537 ( .I1(n15629), .I2(n15628), .I3(n15627), .O(n15638) );
  AOI22S U18538 ( .A1(n20032), .A2(img[567]), .B1(n15630), .B2(img[1591]), .O(
        n15636) );
  MOAI1S U18539 ( .A1(n15668), .A2(n30060), .B1(n13879), .B2(img[439]), .O(
        n15633) );
  MOAI1S U18540 ( .A1(n15631), .A2(n30054), .B1(n19642), .B2(img[183]), .O(
        n15632) );
  NR2 U18541 ( .I1(n15633), .I2(n15632), .O(n15635) );
  AOI22S U18542 ( .A1(n18922), .A2(img[1207]), .B1(n14392), .B2(img[1335]), 
        .O(n15634) );
  ND3S U18543 ( .I1(n15636), .I2(n15635), .I3(n15634), .O(n15637) );
  NR2 U18544 ( .I1(n15638), .I2(n15637), .O(n15827) );
  AOI22S U18545 ( .A1(n15653), .A2(img[1015]), .B1(n19642), .B2(img[247]), .O(
        n15642) );
  AOI22S U18546 ( .A1(n15799), .A2(img[503]), .B1(n15786), .B2(img[375]), .O(
        n15641) );
  AOI22S U18547 ( .A1(n15800), .A2(img[1271]), .B1(n17088), .B2(img[1399]), 
        .O(n15640) );
  AOI22S U18548 ( .A1(n13841), .A2(img[119]), .B1(n13876), .B2(img[631]), .O(
        n15639) );
  MOAI1S U18549 ( .A1(n13850), .A2(n30090), .B1(n20033), .B2(img[2039]), .O(
        n15644) );
  MOAI1S U18550 ( .A1(n15765), .A2(n30078), .B1(n13797), .B2(img[759]), .O(
        n15643) );
  NR2 U18551 ( .I1(n15644), .I2(n15643), .O(n15648) );
  MOAI1S U18552 ( .A1(n15698), .A2(n30086), .B1(n15751), .B2(img[1911]), .O(
        n15646) );
  MOAI1S U18553 ( .A1(n15780), .A2(n30059), .B1(n13885), .B2(img[887]), .O(
        n15645) );
  NR2 U18554 ( .I1(n15646), .I2(n15645), .O(n15647) );
  MOAI1 U18555 ( .A1(n15827), .A2(n15142), .B1(n16236), .B2(n13846), .O(n15707) );
  NR2 U18556 ( .I1(n15651), .I2(n15650), .O(n15656) );
  AOI22S U18557 ( .A1(n13837), .A2(img[687]), .B1(n15652), .B2(img[1711]), .O(
        n15655) );
  AOI22S U18558 ( .A1(n22928), .A2(img[1967]), .B1(n14112), .B2(img[943]), .O(
        n15654) );
  ND3S U18559 ( .I1(n15656), .I2(n15655), .I3(n15654), .O(n15665) );
  MOAI1S U18560 ( .A1(n15698), .A2(n30081), .B1(n15800), .B2(img[1199]), .O(
        n15659) );
  MOAI1S U18561 ( .A1(n15674), .A2(n30228), .B1(n15657), .B2(img[559]), .O(
        n15658) );
  NR2 U18562 ( .I1(n15659), .I2(n15658), .O(n15663) );
  AOI22S U18563 ( .A1(n15799), .A2(img[431]), .B1(n15786), .B2(img[303]), .O(
        n15662) );
  AOI22S U18564 ( .A1(n15660), .A2(img[175]), .B1(n13854), .B2(img[1327]), .O(
        n15661) );
  ND3S U18565 ( .I1(n15663), .I2(n15662), .I3(n15661), .O(n15664) );
  MOAI1S U18566 ( .A1(n13850), .A2(n30222), .B1(n15080), .B2(img[2007]), .O(
        n15671) );
  MOAI1S U18567 ( .A1(n15765), .A2(n30074), .B1(n13797), .B2(img[727]), .O(
        n15670) );
  AOI22S U18568 ( .A1(n13882), .A2(img[471]), .B1(n17880), .B2(img[343]), .O(
        n15667) );
  ND2S U18569 ( .I1(n13885), .I2(img[855]), .O(n15666) );
  OAI112HS U18570 ( .C1(n15668), .C2(n30215), .A1(n15667), .B1(n15666), .O(
        n15669) );
  NR3 U18571 ( .I1(n15671), .I2(n15670), .I3(n15669), .O(n15679) );
  MOAI1S U18572 ( .A1(n13838), .A2(n30199), .B1(n17088), .B2(img[1367]), .O(
        n15673) );
  MOAI1S U18573 ( .A1(n19648), .A2(n30238), .B1(n19642), .B2(img[215]), .O(
        n15672) );
  NR2 U18574 ( .I1(n15673), .I2(n15672), .O(n15678) );
  MOAI1S U18575 ( .A1(n15698), .A2(n30082), .B1(n15751), .B2(img[1879]), .O(
        n15676) );
  MOAI1S U18576 ( .A1(n15674), .A2(n30227), .B1(n13883), .B2(img[599]), .O(
        n15675) );
  NR2 U18577 ( .I1(n15676), .I2(n15675), .O(n15677) );
  ND3 U18578 ( .I1(n15679), .I2(n15678), .I3(n15677), .O(n16227) );
  AOI22S U18579 ( .A1(n15653), .A2(img[935]), .B1(n19642), .B2(img[167]), .O(
        n15683) );
  AOI22S U18580 ( .A1(n15799), .A2(img[423]), .B1(n15786), .B2(img[295]), .O(
        n15682) );
  AOI22S U18581 ( .A1(n15800), .A2(img[1191]), .B1(n14392), .B2(img[1319]), 
        .O(n15681) );
  AOI22S U18582 ( .A1(n18958), .A2(img[39]), .B1(n15657), .B2(img[551]), .O(
        n15680) );
  MOAI1S U18583 ( .A1(n13850), .A2(n30152), .B1(n17514), .B2(img[1959]), .O(
        n15685) );
  MOAI1S U18584 ( .A1(n15765), .A2(n30140), .B1(n13898), .B2(img[679]), .O(
        n15684) );
  NR2 U18585 ( .I1(n15685), .I2(n15684), .O(n15689) );
  MOAI1S U18586 ( .A1(n15698), .A2(n30148), .B1(n15751), .B2(img[1831]), .O(
        n15687) );
  NR2 U18587 ( .I1(n15687), .I2(n15686), .O(n15688) );
  AOI22S U18588 ( .A1(n16227), .A2(n17938), .B1(n16244), .B2(n20124), .O(
        n15705) );
  AOI22S U18589 ( .A1(n15653), .A2(img[1007]), .B1(n19642), .B2(img[239]), .O(
        n15695) );
  AOI22S U18590 ( .A1(n15691), .A2(img[495]), .B1(n17880), .B2(img[367]), .O(
        n15694) );
  AOI22S U18591 ( .A1(n15800), .A2(img[1263]), .B1(n17088), .B2(img[1391]), 
        .O(n15693) );
  AOI22S U18592 ( .A1(n13803), .A2(img[111]), .B1(n15657), .B2(img[623]), .O(
        n15692) );
  MOAI1S U18593 ( .A1(n13850), .A2(n30223), .B1(n15080), .B2(img[2031]), .O(
        n15697) );
  MOAI1S U18594 ( .A1(n15765), .A2(n30076), .B1(n13837), .B2(img[751]), .O(
        n15696) );
  NR2 U18595 ( .I1(n15697), .I2(n15696), .O(n15702) );
  MOAI1S U18596 ( .A1(n15698), .A2(n30084), .B1(n15751), .B2(img[1903]), .O(
        n15700) );
  MOAI1S U18597 ( .A1(n15780), .A2(n30216), .B1(n13885), .B2(img[879]), .O(
        n15699) );
  NR2 U18598 ( .I1(n15700), .I2(n15699), .O(n15701) );
  ND2S U18599 ( .I1(n16246), .I2(n13839), .O(n15704) );
  OAI112HS U18600 ( .C1(n16228), .C2(n16468), .A1(n15705), .B1(n15704), .O(
        n15706) );
  MOAI1S U18601 ( .A1(n19648), .A2(n30207), .B1(n19642), .B2(img[151]), .O(
        n15709) );
  NR2 U18602 ( .I1(n15710), .I2(n15709), .O(n15713) );
  AOI22S U18603 ( .A1(n15800), .A2(img[1175]), .B1(n17088), .B2(img[1303]), 
        .O(n15712) );
  AOI22S U18604 ( .A1(n17778), .A2(img[23]), .B1(n15506), .B2(img[535]), .O(
        n15711) );
  AOI22S U18605 ( .A1(n18885), .A2(img[1815]), .B1(n15630), .B2(img[1559]), 
        .O(n15718) );
  MOAI1S U18606 ( .A1(n13850), .A2(n30224), .B1(n22928), .B2(img[1943]), .O(
        n15715) );
  MOAI1S U18607 ( .A1(n15765), .A2(n30075), .B1(n13797), .B2(img[663]), .O(
        n15714) );
  NR2 U18608 ( .I1(n15715), .I2(n15714), .O(n15717) );
  AOI22S U18609 ( .A1(n13884), .A2(img[791]), .B1(n13845), .B2(img[1431]), .O(
        n15716) );
  ND3S U18610 ( .I1(n15718), .I2(n15717), .I3(n15716), .O(n15719) );
  AOI22S U18611 ( .A1(n15653), .A2(img[999]), .B1(n19642), .B2(img[231]), .O(
        n15725) );
  AOI22S U18612 ( .A1(n13882), .A2(img[487]), .B1(n15786), .B2(img[359]), .O(
        n15724) );
  AOI22S U18613 ( .A1(n15800), .A2(img[1255]), .B1(n17088), .B2(img[1383]), 
        .O(n15723) );
  AOI22S U18614 ( .A1(n18983), .A2(img[103]), .B1(n13876), .B2(img[615]), .O(
        n15722) );
  MOAI1S U18615 ( .A1(n13850), .A2(n30154), .B1(n20033), .B2(img[2023]), .O(
        n15727) );
  MOAI1S U18616 ( .A1(n15765), .A2(n30142), .B1(n13837), .B2(img[743]), .O(
        n15726) );
  NR2 U18617 ( .I1(n15727), .I2(n15726), .O(n15731) );
  NR2 U18618 ( .I1(n15729), .I2(n15728), .O(n15730) );
  MOAI1 U18619 ( .A1(n16239), .A2(n17656), .B1(n16247), .B2(n21062), .O(n15759) );
  MOAI1S U18620 ( .A1(n19648), .A2(n30257), .B1(n19642), .B2(img[143]), .O(
        n15733) );
  AOI22S U18621 ( .A1(n15800), .A2(img[1167]), .B1(n17088), .B2(img[1295]), 
        .O(n15736) );
  AOI22S U18622 ( .A1(n19290), .A2(img[15]), .B1(n20032), .B2(img[527]), .O(
        n15735) );
  AOI22S U18623 ( .A1(n16075), .A2(img[1807]), .B1(n13823), .B2(img[1551]), 
        .O(n15742) );
  MOAI1S U18624 ( .A1(n13850), .A2(n30089), .B1(n20033), .B2(img[1935]), .O(
        n15739) );
  MOAI1S U18625 ( .A1(n15765), .A2(n30077), .B1(n13837), .B2(img[655]), .O(
        n15738) );
  NR2 U18626 ( .I1(n15739), .I2(n15738), .O(n15741) );
  AOI22S U18627 ( .A1(n13884), .A2(img[783]), .B1(n13845), .B2(img[1423]), .O(
        n15740) );
  AOI22S U18628 ( .A1(n15653), .A2(img[967]), .B1(n19642), .B2(img[199]), .O(
        n15748) );
  AOI22S U18629 ( .A1(n15799), .A2(img[455]), .B1(n15786), .B2(img[327]), .O(
        n15747) );
  AOI22S U18630 ( .A1(n15800), .A2(img[1223]), .B1(n14392), .B2(img[1351]), 
        .O(n15746) );
  AOI22S U18631 ( .A1(n17886), .A2(img[71]), .B1(n13876), .B2(img[583]), .O(
        n15745) );
  AN4S U18632 ( .I1(n15748), .I2(n15747), .I3(n15746), .I4(n15745), .O(n15757)
         );
  MOAI1S U18633 ( .A1(n13850), .A2(n30193), .B1(n15080), .B2(img[1991]), .O(
        n15750) );
  MOAI1S U18634 ( .A1(n15806), .A2(n30137), .B1(n13797), .B2(img[711]), .O(
        n15749) );
  NR2 U18635 ( .I1(n15750), .I2(n15749), .O(n15756) );
  MOAI1S U18636 ( .A1(n15698), .A2(n30145), .B1(n15751), .B2(img[1863]), .O(
        n15754) );
  MOAI1S U18637 ( .A1(n15780), .A2(n30187), .B1(n13885), .B2(img[839]), .O(
        n15753) );
  NR2 U18638 ( .I1(n15754), .I2(n15753), .O(n15755) );
  ND3 U18639 ( .I1(n15757), .I2(n15756), .I3(n15755), .O(n16238) );
  MOAI1S U18640 ( .A1(n16241), .A2(n13945), .B1(n16238), .B2(n18040), .O(
        n15758) );
  MOAI1S U18641 ( .A1(n19648), .A2(n30114), .B1(n19642), .B2(img[159]), .O(
        n15760) );
  AOI22S U18642 ( .A1(n15800), .A2(img[1183]), .B1(n14392), .B2(img[1311]), 
        .O(n15763) );
  AOI22S U18643 ( .A1(n17778), .A2(img[31]), .B1(n13876), .B2(img[543]), .O(
        n15762) );
  ND3 U18644 ( .I1(n15764), .I2(n15763), .I3(n15762), .O(n15772) );
  AOI22S U18645 ( .A1(n20038), .A2(img[1823]), .B1(n13823), .B2(img[1567]), 
        .O(n15770) );
  MOAI1S U18646 ( .A1(n13850), .A2(n30155), .B1(n15080), .B2(img[1951]), .O(
        n15767) );
  MOAI1S U18647 ( .A1(n15765), .A2(n30143), .B1(n13797), .B2(img[671]), .O(
        n15766) );
  NR2 U18648 ( .I1(n15767), .I2(n15766), .O(n15769) );
  AOI22S U18649 ( .A1(n19641), .A2(img[799]), .B1(n13845), .B2(img[1439]), .O(
        n15768) );
  ND3S U18650 ( .I1(n15770), .I2(n15769), .I3(n15768), .O(n15771) );
  AOI22S U18651 ( .A1(n15653), .A2(img[1023]), .B1(n15773), .B2(img[255]), .O(
        n15777) );
  AOI22S U18652 ( .A1(n15799), .A2(img[511]), .B1(n13800), .B2(img[383]), .O(
        n15776) );
  AOI22S U18653 ( .A1(n15800), .A2(img[1279]), .B1(n14392), .B2(img[1407]), 
        .O(n15775) );
  AOI22S U18654 ( .A1(n17886), .A2(img[127]), .B1(n13876), .B2(img[639]), .O(
        n15774) );
  MOAI1S U18655 ( .A1(n13850), .A2(n30191), .B1(n22928), .B2(img[2047]), .O(
        n15779) );
  MOAI1S U18656 ( .A1(n15806), .A2(n30139), .B1(n13837), .B2(img[767]), .O(
        n15778) );
  NR2 U18657 ( .I1(n15779), .I2(n15778), .O(n15784) );
  MOAI1S U18658 ( .A1(n15698), .A2(n30147), .B1(n15809), .B2(img[1919]), .O(
        n15782) );
  MOAI1S U18659 ( .A1(n15780), .A2(n30185), .B1(n13886), .B2(img[895]), .O(
        n15781) );
  NR2 U18660 ( .I1(n15782), .I2(n15781), .O(n15783) );
  MOAI1 U18661 ( .A1(n16233), .A2(n13766), .B1(n16245), .B2(n20969), .O(n15816) );
  MOAI1S U18662 ( .A1(n19648), .A2(n30176), .B1(n19642), .B2(img[191]), .O(
        n15787) );
  NR2 U18663 ( .I1(n15788), .I2(n15787), .O(n15791) );
  AOI22S U18664 ( .A1(n13787), .A2(img[1215]), .B1(n16799), .B2(img[1343]), 
        .O(n15790) );
  AOI22S U18665 ( .A1(n17864), .A2(img[63]), .B1(n13876), .B2(img[575]), .O(
        n15789) );
  ND3 U18666 ( .I1(n15791), .I2(n15790), .I3(n15789), .O(n15798) );
  AOI22S U18667 ( .A1(n13870), .A2(img[1855]), .B1(n18837), .B2(img[1599]), 
        .O(n15796) );
  MOAI1S U18668 ( .A1(n13850), .A2(n30192), .B1(n17514), .B2(img[1983]), .O(
        n15793) );
  MOAI1S U18669 ( .A1(n15806), .A2(n30136), .B1(n13837), .B2(img[703]), .O(
        n15792) );
  NR2 U18670 ( .I1(n15793), .I2(n15792), .O(n15795) );
  AOI22S U18671 ( .A1(n15568), .A2(img[831]), .B1(n13845), .B2(img[1471]), .O(
        n15794) );
  ND3S U18672 ( .I1(n15796), .I2(n15795), .I3(n15794), .O(n15797) );
  AOI22S U18673 ( .A1(n15653), .A2(img[975]), .B1(n19642), .B2(img[207]), .O(
        n15805) );
  AOI22S U18674 ( .A1(n15799), .A2(img[463]), .B1(n19710), .B2(img[335]), .O(
        n15804) );
  AOI22S U18675 ( .A1(n15800), .A2(img[1231]), .B1(n17088), .B2(img[1359]), 
        .O(n15803) );
  AOI22S U18676 ( .A1(n13803), .A2(img[79]), .B1(n13876), .B2(img[591]), .O(
        n15802) );
  MOAI1S U18677 ( .A1(n13850), .A2(n30092), .B1(n15080), .B2(img[1999]), .O(
        n15808) );
  MOAI1S U18678 ( .A1(n15806), .A2(n30080), .B1(n13898), .B2(img[719]), .O(
        n15807) );
  NR2 U18679 ( .I1(n15808), .I2(n15807), .O(n15813) );
  MOAI1S U18680 ( .A1(n15698), .A2(n30088), .B1(n15809), .B2(img[1871]), .O(
        n15811) );
  MOAI1S U18681 ( .A1(n15780), .A2(n30061), .B1(n13885), .B2(img[847]), .O(
        n15810) );
  NR2 U18682 ( .I1(n15811), .I2(n15810), .O(n15812) );
  MOAI1 U18683 ( .A1(n15828), .A2(n17658), .B1(n16234), .B2(n20263), .O(n15815) );
  NR2 U18684 ( .I1(n15816), .I2(n15815), .O(n15817) );
  NR2 U18685 ( .I1(n17656), .I2(n16233), .O(n15821) );
  NR2 U18686 ( .I1(n15821), .I2(n15820), .O(n15824) );
  AOI22S U18687 ( .A1(n16245), .A2(n13846), .B1(n20438), .B2(n16244), .O(
        n15823) );
  AOI22S U18688 ( .A1(n16229), .A2(n17938), .B1(n20406), .B2(n16247), .O(
        n15822) );
  ND3S U18689 ( .I1(n15824), .I2(n15823), .I3(n15822), .O(n15833) );
  MOAI1S U18690 ( .A1(n16239), .A2(n13945), .B1(n16234), .B2(n18040), .O(
        n15825) );
  NR2 U18691 ( .I1(n15826), .I2(n15825), .O(n15831) );
  INV1S U18692 ( .I(n15827), .O(n16237) );
  AOI22S U18693 ( .A1(n13839), .A2(n16236), .B1(n16237), .B2(n17875), .O(
        n15830) );
  INV1S U18694 ( .I(n15828), .O(n16240) );
  INV2 U18695 ( .I(n15142), .O(n20187) );
  AOI22S U18696 ( .A1(n21062), .A2(n16246), .B1(n16240), .B2(n20187), .O(
        n15829) );
  NR2 U18697 ( .I1(n15833), .I2(n15832), .O(n15834) );
  NR2 U18698 ( .I1(n20969), .I2(n15834), .O(n19452) );
  NR2 U18699 ( .I1(n21800), .I2(n21238), .O(n15902) );
  NR2 U18700 ( .I1(n21728), .I2(n15867), .O(n15877) );
  INV1S U18701 ( .I(template_store[47]), .O(n21727) );
  NR2 U18702 ( .I1(n21727), .I2(n21799), .O(n15876) );
  NR2 U18703 ( .I1(n15868), .I2(n21231), .O(n15891) );
  NR2 U18704 ( .I1(n21730), .I2(n15886), .O(n15890) );
  FA1 U18705 ( .A(n15845), .B(n15844), .CI(n15843), .CO(n21778), .S(n21780) );
  NR2 U18706 ( .I1(n15878), .I2(n15886), .O(n15855) );
  NR2 U18707 ( .I1(n21800), .I2(n15867), .O(n15852) );
  NR2 U18708 ( .I1(n15878), .I2(n21799), .O(n15851) );
  NR2 U18709 ( .I1(n15875), .I2(n15867), .O(n15847) );
  NR2 U18710 ( .I1(n15868), .I2(n21799), .O(n15846) );
  NR2 U18711 ( .I1(n15875), .I2(n21336), .O(n15857) );
  FA1 U18712 ( .A(n15850), .B(n15849), .CI(n15848), .CO(n15860), .S(n15856) );
  NR2 U18713 ( .I1(n21800), .I2(n21336), .O(n21787) );
  NR2 U18714 ( .I1(n15875), .I2(n15886), .O(n21790) );
  NR2 U18715 ( .I1(n15875), .I2(n21799), .O(n21792) );
  NR2 U18716 ( .I1(n21800), .I2(n15886), .O(n21791) );
  INV1S U18717 ( .I(n15920), .O(n15863) );
  NR2 U18718 ( .I1(n15918), .I2(n15917), .O(n15862) );
  MOAI1 U18719 ( .A1(n15863), .A2(n15862), .B1(n15917), .B2(n15918), .O(n21779) );
  NR2 U18720 ( .I1(n15885), .I2(n21729), .O(n15871) );
  NR2 U18721 ( .I1(n21727), .I2(n21336), .O(n15870) );
  NR2 U18722 ( .I1(n21728), .I2(n21726), .O(n15866) );
  NR2 U18723 ( .I1(n21730), .I2(n21231), .O(n15865) );
  NR2 U18724 ( .I1(n15868), .I2(n21238), .O(n15864) );
  NR2 U18725 ( .I1(n21728), .I2(n21729), .O(n21742) );
  FA1S U18726 ( .A(n15866), .B(n15865), .CI(n15864), .CO(n21741), .S(n15869)
         );
  NR2 U18727 ( .I1(n21730), .I2(n21726), .O(n21736) );
  NR2 U18728 ( .I1(n21727), .I2(n21231), .O(n21735) );
  NR2 U18729 ( .I1(n15885), .I2(n21238), .O(n21734) );
  NR2 U18730 ( .I1(n21727), .I2(n15867), .O(n15874) );
  NR2 U18731 ( .I1(n15878), .I2(n21238), .O(n15873) );
  NR2 U18732 ( .I1(n21730), .I2(n15867), .O(n15888) );
  NR2 U18733 ( .I1(n15885), .I2(n21726), .O(n15884) );
  NR2 U18734 ( .I1(n21728), .I2(n21231), .O(n15883) );
  NR2 U18735 ( .I1(n15868), .I2(n21729), .O(n15882) );
  FA1S U18736 ( .A(n15871), .B(n15870), .CI(n15869), .CO(n21748), .S(n15879)
         );
  NR2 U18737 ( .I1(n21730), .I2(n21336), .O(n15897) );
  NR2 U18738 ( .I1(n15875), .I2(n21238), .O(n15894) );
  NR2 U18739 ( .I1(n15878), .I2(n21729), .O(n15892) );
  FA1S U18740 ( .A(n15881), .B(n15880), .CI(n15879), .CO(n21746), .S(n15911)
         );
  NR2 U18741 ( .I1(n15885), .I2(n21231), .O(n15900) );
  NR2 U18742 ( .I1(n21727), .I2(n15886), .O(n15899) );
  HA1 U18743 ( .A(n15888), .B(n15887), .C(n15872), .S(n15898) );
  NR2 U18744 ( .I1(n21728), .I2(n21336), .O(n21766) );
  XNR2HS U18745 ( .I1(n21750), .I2(n21751), .O(n15916) );
  FA1 U18746 ( .A(n15897), .B(n15896), .CI(n15895), .CO(n15912), .S(n21795) );
  FA1 U18747 ( .A(n15906), .B(n15905), .CI(n15904), .CO(n21770), .S(n21775) );
  FA1 U18748 ( .A(n15909), .B(n15908), .CI(n15907), .CO(n15910), .S(n21793) );
  FA1S U18749 ( .A(n15912), .B(n15911), .CI(n15910), .CO(n21751), .S(n21631)
         );
  AOI12H U18750 ( .B1(mult_x_431_n11), .B2(mult_x_431_n7), .A1(n15914), .O(
        n21634) );
  MOAI1H U18751 ( .A1(n15915), .A2(n21634), .B1(n21632), .B2(n21631), .O(
        n21749) );
  XNR2HS U18752 ( .I1(n15916), .I2(n21749), .O(PE_N59) );
  XNR2HS U18753 ( .I1(n15918), .I2(n15917), .O(n15919) );
  XNR2HS U18754 ( .I1(n15920), .I2(n15919), .O(PE_N53) );
  INV1S U18755 ( .I(template_store[34]), .O(n15979) );
  INV1S U18756 ( .I(n21254), .O(n23525) );
  NR2 U18757 ( .I1(n15979), .I2(n23525), .O(n15930) );
  INV1S U18758 ( .I(n21259), .O(n23537) );
  INV1S U18759 ( .I(template_store[33]), .O(n15986) );
  NR2 U18760 ( .I1(n23537), .I2(n15986), .O(n15929) );
  INV1S U18761 ( .I(template_store[39]), .O(n23536) );
  NR2 U18762 ( .I1(n23536), .I2(n22942), .O(n15926) );
  NR2 U18763 ( .I1(n15979), .I2(n23508), .O(n15925) );
  INV1S U18764 ( .I(template_store[38]), .O(n23526) );
  NR2 U18765 ( .I1(n23526), .I2(n15985), .O(n15924) );
  INV1S U18766 ( .I(template_store[37]), .O(n23509) );
  NR2 U18767 ( .I1(n23509), .I2(n13818), .O(n15923) );
  INV1S U18768 ( .I(template_store[35]), .O(n23480) );
  NR2 U18769 ( .I1(n23480), .I2(n13817), .O(n15922) );
  INV1S U18770 ( .I(template_store[36]), .O(n23490) );
  NR2 U18771 ( .I1(n23490), .I2(n13816), .O(n15921) );
  FA1S U18772 ( .A(n15923), .B(n15922), .CI(n15921), .CO(n15940), .S(n15953)
         );
  NR2 U18773 ( .I1(n23490), .I2(n13818), .O(n15967) );
  NR2 U18774 ( .I1(n23480), .I2(n13816), .O(n15966) );
  NR2 U18775 ( .I1(n15986), .I2(n13817), .O(n15961) );
  INV1S U18776 ( .I(template_store[32]), .O(n23470) );
  NR2 U18777 ( .I1(n23470), .I2(n23508), .O(n15960) );
  NR2 U18778 ( .I1(n23490), .I2(n13817), .O(n15933) );
  NR2 U18779 ( .I1(n23480), .I2(n23508), .O(n15932) );
  NR2 U18780 ( .I1(n23536), .I2(n15985), .O(n15931) );
  NR2 U18781 ( .I1(n23526), .I2(n13818), .O(n15939) );
  NR2 U18782 ( .I1(n23509), .I2(n13816), .O(n15938) );
  NR2 U18783 ( .I1(n23537), .I2(n23470), .O(n15927) );
  NR2 U18784 ( .I1(n15986), .I2(n23508), .O(n15944) );
  NR2 U18785 ( .I1(n23470), .I2(n23525), .O(n15943) );
  HA1 U18786 ( .A(n15928), .B(n15927), .C(n15937), .S(n15949) );
  NR2 U18787 ( .I1(n23526), .I2(n22942), .O(n15947) );
  NR2 U18788 ( .I1(n15979), .I2(n13817), .O(n15946) );
  NR2 U18789 ( .I1(n23509), .I2(n15985), .O(n15945) );
  HA1 U18790 ( .A(n15930), .B(n15929), .C(n23483), .S(n15942) );
  FA1S U18791 ( .A(n15933), .B(n15932), .CI(n15931), .CO(n23482), .S(n15936)
         );
  NR2 U18792 ( .I1(n23490), .I2(n23508), .O(n23479) );
  NR2 U18793 ( .I1(n23509), .I2(n13817), .O(n23478) );
  NR2 U18794 ( .I1(n23526), .I2(n13816), .O(n23477) );
  FA1S U18795 ( .A(n15936), .B(n15935), .CI(n15934), .CO(n23495), .S(n15954)
         );
  NR2 U18796 ( .I1(n23536), .I2(n13818), .O(n23473) );
  NR2 U18797 ( .I1(n23537), .I2(n15979), .O(n23472) );
  NR2 U18798 ( .I1(n23480), .I2(n23525), .O(n23471) );
  FA1S U18799 ( .A(n15939), .B(n15938), .CI(n15937), .CO(n23475), .S(n15935)
         );
  FA1S U18800 ( .A(n15942), .B(n15941), .CI(n15940), .CO(n23474), .S(n15956)
         );
  XNR2HS U18801 ( .I1(n23501), .I2(n23502), .O(n16000) );
  HA1 U18802 ( .A(n15944), .B(n15943), .C(n15950), .S(n15970) );
  NR2 U18803 ( .I1(n23509), .I2(n22942), .O(n15959) );
  NR2 U18804 ( .I1(n15979), .I2(n13816), .O(n15958) );
  NR2 U18805 ( .I1(n23480), .I2(n13818), .O(n15957) );
  FA1S U18806 ( .A(n15947), .B(n15946), .CI(n15945), .CO(n15948), .S(n15968)
         );
  FA1S U18807 ( .A(n15950), .B(n15949), .CI(n15948), .CO(n15934), .S(n15996)
         );
  FA1S U18808 ( .A(n15956), .B(n15955), .CI(n15954), .CO(n23501), .S(n23523)
         );
  NR2 U18809 ( .I1(n23490), .I2(n22942), .O(n15975) );
  NR2 U18810 ( .I1(n15979), .I2(n13818), .O(n15974) );
  NR2 U18811 ( .I1(n23480), .I2(n15985), .O(n15973) );
  FA1S U18812 ( .A(n15959), .B(n15958), .CI(n15957), .CO(n15969), .S(n15977)
         );
  NR2 U18813 ( .I1(n23490), .I2(n15985), .O(n15964) );
  NR2 U18814 ( .I1(n15986), .I2(n13816), .O(n15972) );
  NR2 U18815 ( .I1(n23470), .I2(n13817), .O(n15971) );
  FA1S U18816 ( .A(n15967), .B(n15966), .CI(n15965), .CO(n15951), .S(n15993)
         );
  FA1S U18817 ( .A(n15970), .B(n15969), .CI(n15968), .CO(n15997), .S(n15992)
         );
  NR2 U18818 ( .I1(n15986), .I2(n13818), .O(n15984) );
  NR2 U18819 ( .I1(n23470), .I2(n13816), .O(n15983) );
  HA1 U18820 ( .A(n15972), .B(n15971), .C(n15963), .S(n15981) );
  FA1S U18821 ( .A(n15975), .B(n15974), .CI(n15973), .CO(n15978), .S(n15980)
         );
  FA1 U18822 ( .A(n15978), .B(n15977), .CI(n15976), .CO(n23552), .S(n23548) );
  NR2 U18823 ( .I1(n23480), .I2(n22942), .O(n15991) );
  NR2 U18824 ( .I1(n15979), .I2(n15985), .O(n15990) );
  NR2 U18825 ( .I1(n15979), .I2(n22942), .O(n15988) );
  NR2 U18826 ( .I1(n15986), .I2(n15985), .O(n15987) );
  FA1 U18827 ( .A(n15982), .B(n15981), .CI(n15980), .CO(n23549), .S(n23557) );
  NR2 U18828 ( .I1(n23470), .I2(n13818), .O(n23555) );
  NR2 U18829 ( .I1(n23470), .I2(n15985), .O(n23469) );
  NR2 U18830 ( .I1(n15986), .I2(n22942), .O(n23468) );
  FA1S U18831 ( .A(n15991), .B(n15990), .CI(n15989), .CO(n23558), .S(n21723)
         );
  INV1S U18832 ( .I(n21630), .O(n15999) );
  FA1 U18833 ( .A(n15994), .B(n15993), .CI(n15992), .CO(n21628), .S(n23551) );
  FA1S U18834 ( .A(n15997), .B(n15996), .CI(n15995), .CO(n23524), .S(n21627)
         );
  NR2 U18835 ( .I1(n21628), .I2(n21627), .O(n15998) );
  MOAI1 U18836 ( .A1(n15999), .A2(n15998), .B1(n21627), .B2(n21628), .O(n23522) );
  XNR2HS U18837 ( .I1(n16000), .I2(n23500), .O(PE_N73) );
  AOI22S U18838 ( .A1(n18681), .A2(img[495]), .B1(n13855), .B2(img[367]), .O(
        n16007) );
  AOI22S U18839 ( .A1(n18935), .A2(img[1007]), .B1(n13893), .B2(img[879]), .O(
        n16006) );
  BUF1 U18840 ( .I(n13800), .O(n17377) );
  AOI22S U18841 ( .A1(n17377), .A2(img[239]), .B1(n17376), .B2(img[111]), .O(
        n16005) );
  AOI22S U18842 ( .A1(n19641), .A2(img[751]), .B1(n13797), .B2(img[623]), .O(
        n16004) );
  AN4S U18843 ( .I1(n16007), .I2(n16006), .I3(n16005), .I4(n16004), .O(n16015)
         );
  AOI22S U18844 ( .A1(n17382), .A2(img[1519]), .B1(n13845), .B2(img[1391]), 
        .O(n16013) );
  BUF6 U18845 ( .I(n20033), .O(n17383) );
  AOI22S U18846 ( .A1(n17864), .A2(img[2031]), .B1(n17383), .B2(img[1903]), 
        .O(n16012) );
  INV1S U18847 ( .I(n13789), .O(n17323) );
  AOI22S U18848 ( .A1(n17323), .A2(img[1263]), .B1(n18974), .B2(img[1135]), 
        .O(n16011) );
  AOI22S U18849 ( .A1(n19036), .A2(img[1775]), .B1(n13794), .B2(img[1647]), 
        .O(n16010) );
  AN4S U18850 ( .I1(n16013), .I2(n16012), .I3(n16011), .I4(n16010), .O(n16014)
         );
  AOI22S U18851 ( .A1(n20102), .A2(img[431]), .B1(n13858), .B2(img[303]), .O(
        n16020) );
  AOI22S U18852 ( .A1(n19037), .A2(img[943]), .B1(n13890), .B2(img[815]), .O(
        n16019) );
  BUF1 U18853 ( .I(n13800), .O(n17271) );
  AOI22S U18854 ( .A1(n17271), .A2(img[175]), .B1(n17376), .B2(img[47]), .O(
        n16018) );
  AOI22S U18855 ( .A1(n16348), .A2(img[687]), .B1(n13898), .B2(img[559]), .O(
        n16017) );
  AN4S U18856 ( .I1(n16020), .I2(n16019), .I3(n16018), .I4(n16017), .O(n16026)
         );
  AOI22S U18857 ( .A1(n19193), .A2(img[1455]), .B1(n16127), .B2(img[1327]), 
        .O(n16024) );
  AOI22S U18858 ( .A1(n13833), .A2(img[1967]), .B1(n17383), .B2(img[1839]), 
        .O(n16023) );
  INV1S U18859 ( .I(n13789), .O(n17277) );
  AOI22S U18860 ( .A1(n17277), .A2(img[1199]), .B1(n17276), .B2(img[1071]), 
        .O(n16022) );
  AOI22S U18861 ( .A1(n19215), .A2(img[1711]), .B1(n13794), .B2(img[1583]), 
        .O(n16021) );
  AN4S U18862 ( .I1(n16024), .I2(n16023), .I3(n16022), .I4(n16021), .O(n16025)
         );
  AOI22S U18863 ( .A1(n20611), .A2(n13839), .B1(n17875), .B2(n20610), .O(
        n16092) );
  AOI22S U18864 ( .A1(n13785), .A2(img[439]), .B1(n13858), .B2(img[311]), .O(
        n16030) );
  AOI22S U18865 ( .A1(n18148), .A2(img[951]), .B1(n13890), .B2(img[823]), .O(
        n16029) );
  AOI22S U18866 ( .A1(n18818), .A2(img[183]), .B1(n17376), .B2(img[55]), .O(
        n16028) );
  AOI22S U18867 ( .A1(n13826), .A2(img[695]), .B1(n13837), .B2(img[567]), .O(
        n16027) );
  AN4S U18868 ( .I1(n16030), .I2(n16029), .I3(n16028), .I4(n16027), .O(n16036)
         );
  AOI22S U18869 ( .A1(n15630), .A2(img[1463]), .B1(n17827), .B2(img[1335]), 
        .O(n16034) );
  AOI22S U18870 ( .A1(n17864), .A2(img[1975]), .B1(n17383), .B2(img[1847]), 
        .O(n16033) );
  AOI22S U18871 ( .A1(n16635), .A2(img[1207]), .B1(n19647), .B2(img[1079]), 
        .O(n16032) );
  AOI22S U18872 ( .A1(n19215), .A2(img[1719]), .B1(n17550), .B2(img[1591]), 
        .O(n16031) );
  AN4S U18873 ( .I1(n16034), .I2(n16033), .I3(n16032), .I4(n16031), .O(n16035)
         );
  AOI22S U18874 ( .A1(n20102), .A2(img[487]), .B1(n13855), .B2(img[359]), .O(
        n16041) );
  AOI22S U18875 ( .A1(n19956), .A2(img[999]), .B1(n17115), .B2(img[871]), .O(
        n16040) );
  BUF1 U18876 ( .I(n13800), .O(n17197) );
  AOI22S U18877 ( .A1(n17197), .A2(img[231]), .B1(n17376), .B2(img[103]), .O(
        n16039) );
  AOI22S U18878 ( .A1(n19252), .A2(img[743]), .B1(n13797), .B2(img[615]), .O(
        n16038) );
  AN4S U18879 ( .I1(n16041), .I2(n16040), .I3(n16039), .I4(n16038), .O(n16047)
         );
  AOI22S U18880 ( .A1(n19193), .A2(img[1511]), .B1(n19182), .B2(img[1383]), 
        .O(n16045) );
  AOI22S U18881 ( .A1(n17335), .A2(img[2023]), .B1(n17383), .B2(img[1895]), 
        .O(n16044) );
  AOI22S U18882 ( .A1(n18975), .A2(img[1255]), .B1(n15800), .B2(img[1127]), 
        .O(n16043) );
  AOI22S U18883 ( .A1(n19036), .A2(img[1767]), .B1(n13794), .B2(img[1639]), 
        .O(n16042) );
  AN4S U18884 ( .I1(n16045), .I2(n16044), .I3(n16043), .I4(n16042), .O(n16046)
         );
  AOI22S U18885 ( .A1(n20619), .A2(n20187), .B1(n21062), .B2(n20609), .O(
        n16206) );
  AOI22S U18886 ( .A1(n13825), .A2(img[423]), .B1(n13858), .B2(img[295]), .O(
        n16052) );
  AOI22S U18887 ( .A1(n19649), .A2(img[935]), .B1(n16048), .B2(img[807]), .O(
        n16051) );
  AOI22S U18888 ( .A1(n19949), .A2(img[167]), .B1(n17376), .B2(img[39]), .O(
        n16050) );
  AOI22S U18889 ( .A1(n19326), .A2(img[679]), .B1(n13797), .B2(img[551]), .O(
        n16049) );
  AN4S U18890 ( .I1(n16052), .I2(n16051), .I3(n16050), .I4(n16049), .O(n16058)
         );
  AOI22S U18891 ( .A1(n13823), .A2(img[1447]), .B1(n16127), .B2(img[1319]), 
        .O(n16056) );
  AOI22S U18892 ( .A1(n17778), .A2(img[1959]), .B1(n17383), .B2(img[1831]), 
        .O(n16055) );
  AOI22S U18893 ( .A1(n17336), .A2(img[1191]), .B1(n13787), .B2(img[1063]), 
        .O(n16054) );
  AOI22S U18894 ( .A1(n13863), .A2(img[1703]), .B1(n13794), .B2(img[1575]), 
        .O(n16053) );
  AN4S U18895 ( .I1(n16056), .I2(n16055), .I3(n16054), .I4(n16053), .O(n16057)
         );
  ND2 U18896 ( .I1(n16058), .I2(n16057), .O(n20626) );
  AOI22S U18897 ( .A1(n13825), .A2(img[407]), .B1(n13858), .B2(img[279]), .O(
        n16063) );
  AOI22S U18898 ( .A1(n18911), .A2(img[919]), .B1(n13893), .B2(img[791]), .O(
        n16062) );
  BUF1 U18899 ( .I(n13800), .O(n17330) );
  AOI22S U18900 ( .A1(n17330), .A2(img[151]), .B1(n17376), .B2(img[23]), .O(
        n16061) );
  AOI22S U18901 ( .A1(n17835), .A2(img[663]), .B1(n13898), .B2(img[535]), .O(
        n16060) );
  AN4S U18902 ( .I1(n16063), .I2(n16062), .I3(n16061), .I4(n16060), .O(n16070)
         );
  AOI22S U18903 ( .A1(n19193), .A2(img[1431]), .B1(n16127), .B2(img[1303]), 
        .O(n16068) );
  AOI22S U18904 ( .A1(n17793), .A2(img[1943]), .B1(n17383), .B2(img[1815]), 
        .O(n16067) );
  AOI22S U18905 ( .A1(n17336), .A2(img[1175]), .B1(n18922), .B2(img[1047]), 
        .O(n16066) );
  AOI22S U18906 ( .A1(n13863), .A2(img[1687]), .B1(n13794), .B2(img[1559]), 
        .O(n16065) );
  AN4S U18907 ( .I1(n16068), .I2(n16067), .I3(n16066), .I4(n16065), .O(n16069)
         );
  ND2 U18908 ( .I1(n16070), .I2(n16069), .O(n20621) );
  AOI22S U18909 ( .A1(n20626), .A2(n20613), .B1(n17762), .B2(n20621), .O(
        n16208) );
  AOI22S U18910 ( .A1(n13883), .A2(img[399]), .B1(n13858), .B2(img[271]), .O(
        n16074) );
  AOI22S U18911 ( .A1(n16515), .A2(img[911]), .B1(n16048), .B2(img[783]), .O(
        n16073) );
  BUF1 U18912 ( .I(n13800), .O(n17249) );
  AOI22S U18913 ( .A1(n17249), .A2(img[143]), .B1(n17376), .B2(img[15]), .O(
        n16072) );
  AOI22S U18914 ( .A1(n18702), .A2(img[655]), .B1(n13797), .B2(img[527]), .O(
        n16071) );
  AN4S U18915 ( .I1(n16074), .I2(n16073), .I3(n16072), .I4(n16071), .O(n16081)
         );
  AOI22S U18916 ( .A1(n13874), .A2(img[1423]), .B1(n16127), .B2(img[1295]), 
        .O(n16079) );
  AOI22S U18917 ( .A1(n13803), .A2(img[1935]), .B1(n17383), .B2(img[1807]), 
        .O(n16078) );
  INV1S U18918 ( .I(n13789), .O(n18298) );
  AOI22S U18919 ( .A1(n18298), .A2(img[1167]), .B1(n19271), .B2(img[1039]), 
        .O(n16077) );
  AOI22S U18920 ( .A1(n16075), .A2(img[1679]), .B1(n17550), .B2(img[1551]), 
        .O(n16076) );
  AN4S U18921 ( .I1(n16079), .I2(n16078), .I3(n16077), .I4(n16076), .O(n16080)
         );
  ND2 U18922 ( .I1(n16081), .I2(n16080), .O(n20624) );
  AOI22S U18923 ( .A1(n20102), .A2(img[447]), .B1(n13858), .B2(img[319]), .O(
        n16085) );
  AOI22S U18924 ( .A1(n18935), .A2(img[959]), .B1(n13892), .B2(img[831]), .O(
        n16084) );
  AOI22S U18925 ( .A1(n17197), .A2(img[191]), .B1(n17376), .B2(img[63]), .O(
        n16083) );
  AOI22S U18926 ( .A1(n19288), .A2(img[703]), .B1(n13797), .B2(img[575]), .O(
        n16082) );
  AN4S U18927 ( .I1(n16085), .I2(n16084), .I3(n16083), .I4(n16082), .O(n16091)
         );
  AOI22S U18928 ( .A1(n19193), .A2(img[1471]), .B1(n19182), .B2(img[1343]), 
        .O(n16089) );
  AOI22S U18929 ( .A1(n17335), .A2(img[1983]), .B1(n17383), .B2(img[1855]), 
        .O(n16088) );
  INV1S U18930 ( .I(n13789), .O(n17359) );
  AOI22S U18931 ( .A1(n17359), .A2(img[1215]), .B1(n19647), .B2(img[1087]), 
        .O(n16087) );
  AOI22S U18932 ( .A1(n15751), .A2(img[1727]), .B1(n17561), .B2(img[1599]), 
        .O(n16086) );
  AN4S U18933 ( .I1(n16089), .I2(n16088), .I3(n16087), .I4(n16086), .O(n16090)
         );
  ND2 U18934 ( .I1(n16091), .I2(n16090), .O(n20628) );
  AOI22S U18935 ( .A1(n20624), .A2(n13830), .B1(n17928), .B2(n20628), .O(
        n16207) );
  AN4S U18936 ( .I1(n16092), .I2(n16206), .I3(n16208), .I4(n16207), .O(n16168)
         );
  AOI22S U18937 ( .A1(n15506), .A2(img[463]), .B1(n13855), .B2(img[335]), .O(
        n16096) );
  AOI22S U18938 ( .A1(n19956), .A2(img[975]), .B1(n13893), .B2(img[847]), .O(
        n16095) );
  BUF1 U18939 ( .I(n13800), .O(n17354) );
  AOI22S U18940 ( .A1(n17354), .A2(img[207]), .B1(n17376), .B2(img[79]), .O(
        n16094) );
  AOI22S U18941 ( .A1(n19641), .A2(img[719]), .B1(n13898), .B2(img[591]), .O(
        n16093) );
  AN4S U18942 ( .I1(n16096), .I2(n16095), .I3(n16094), .I4(n16093), .O(n16102)
         );
  AOI22S U18943 ( .A1(n17382), .A2(img[1487]), .B1(n18751), .B2(img[1359]), 
        .O(n16100) );
  AOI22S U18944 ( .A1(n17778), .A2(img[1999]), .B1(n17383), .B2(img[1871]), 
        .O(n16099) );
  INV1S U18945 ( .I(n13789), .O(n17347) );
  AOI22S U18946 ( .A1(n17347), .A2(img[1231]), .B1(n13787), .B2(img[1103]), 
        .O(n16098) );
  AOI22S U18947 ( .A1(n15751), .A2(img[1743]), .B1(n18201), .B2(img[1615]), 
        .O(n16097) );
  AN4S U18948 ( .I1(n16100), .I2(n16099), .I3(n16098), .I4(n16097), .O(n16101)
         );
  ND2 U18949 ( .I1(n16102), .I2(n16101), .O(n20614) );
  AOI22S U18950 ( .A1(n13785), .A2(img[391]), .B1(n13858), .B2(img[263]), .O(
        n16106) );
  AOI22S U18951 ( .A1(n14822), .A2(img[903]), .B1(n13890), .B2(img[775]), .O(
        n16105) );
  AOI22S U18952 ( .A1(n17249), .A2(img[135]), .B1(n17376), .B2(img[7]), .O(
        n16104) );
  AOI22S U18953 ( .A1(n16348), .A2(img[647]), .B1(n13837), .B2(img[519]), .O(
        n16103) );
  AN4S U18954 ( .I1(n16106), .I2(n16105), .I3(n16104), .I4(n16103), .O(n16112)
         );
  AOI22S U18955 ( .A1(n17382), .A2(img[1415]), .B1(n16127), .B2(img[1287]), 
        .O(n16110) );
  AOI22S U18956 ( .A1(n13841), .A2(img[1927]), .B1(n17383), .B2(img[1799]), 
        .O(n16109) );
  INV1S U18957 ( .I(n13789), .O(n17254) );
  AOI22S U18958 ( .A1(n17254), .A2(img[1159]), .B1(n19295), .B2(img[1031]), 
        .O(n16108) );
  AOI22S U18959 ( .A1(n19023), .A2(img[1671]), .B1(n13796), .B2(img[1543]), 
        .O(n16107) );
  AN4S U18960 ( .I1(n16110), .I2(n16109), .I3(n16108), .I4(n16107), .O(n16111)
         );
  ND2 U18961 ( .I1(n16112), .I2(n16111), .O(n20627) );
  AOI22S U18962 ( .A1(n20614), .A2(n20263), .B1(n13847), .B2(n20627), .O(
        n16167) );
  AOI22S U18963 ( .A1(n13876), .A2(img[455]), .B1(n13858), .B2(img[327]), .O(
        n16116) );
  AOI22S U18964 ( .A1(n14822), .A2(img[967]), .B1(n13893), .B2(img[839]), .O(
        n16115) );
  AOI22S U18965 ( .A1(n17197), .A2(img[199]), .B1(n17376), .B2(img[71]), .O(
        n16114) );
  AOI22S U18966 ( .A1(n13875), .A2(img[711]), .B1(n13898), .B2(img[583]), .O(
        n16113) );
  AN4S U18967 ( .I1(n16116), .I2(n16115), .I3(n16114), .I4(n16113), .O(n16122)
         );
  AOI22S U18968 ( .A1(n13823), .A2(img[1479]), .B1(n17827), .B2(img[1351]), 
        .O(n16120) );
  AOI22S U18969 ( .A1(n18773), .A2(img[1991]), .B1(n17383), .B2(img[1863]), 
        .O(n16119) );
  AOI22S U18970 ( .A1(n16635), .A2(img[1223]), .B1(n19647), .B2(img[1095]), 
        .O(n16118) );
  AOI22S U18971 ( .A1(n19215), .A2(img[1735]), .B1(n13794), .B2(img[1607]), 
        .O(n16117) );
  AN4S U18972 ( .I1(n16120), .I2(n16119), .I3(n16118), .I4(n16117), .O(n16121)
         );
  ND2 U18973 ( .I1(n16122), .I2(n16121), .O(n20606) );
  BUF1 U18974 ( .I(n18040), .O(n20524) );
  AOI22S U18975 ( .A1(n20102), .A2(img[415]), .B1(n13858), .B2(img[287]), .O(
        n16126) );
  AOI22S U18976 ( .A1(n16037), .A2(img[927]), .B1(n13880), .B2(img[799]), .O(
        n16125) );
  AOI22S U18977 ( .A1(n17788), .A2(img[159]), .B1(n17376), .B2(img[31]), .O(
        n16124) );
  AOI22S U18978 ( .A1(n19641), .A2(img[671]), .B1(n13837), .B2(img[543]), .O(
        n16123) );
  AN4S U18979 ( .I1(n16126), .I2(n16125), .I3(n16124), .I4(n16123), .O(n16133)
         );
  AOI22S U18980 ( .A1(n13823), .A2(img[1439]), .B1(n16127), .B2(img[1311]), 
        .O(n16131) );
  AOI22S U18981 ( .A1(n17515), .A2(img[1951]), .B1(n17383), .B2(img[1823]), 
        .O(n16130) );
  AOI22S U18982 ( .A1(n17277), .A2(img[1183]), .B1(n13787), .B2(img[1055]), 
        .O(n16129) );
  AOI22S U18983 ( .A1(n19215), .A2(img[1695]), .B1(n13794), .B2(img[1567]), 
        .O(n16128) );
  AN4S U18984 ( .I1(n16131), .I2(n16130), .I3(n16129), .I4(n16128), .O(n16132)
         );
  ND2 U18985 ( .I1(n16133), .I2(n16132), .O(n20612) );
  AOI22S U18986 ( .A1(n18681), .A2(img[503]), .B1(n18262), .B2(img[375]), .O(
        n16137) );
  AOI22S U18987 ( .A1(n13788), .A2(img[1015]), .B1(n13893), .B2(img[887]), .O(
        n16136) );
  AOI22S U18988 ( .A1(n19266), .A2(img[247]), .B1(n17376), .B2(img[119]), .O(
        n16135) );
  AOI22S U18989 ( .A1(n16348), .A2(img[759]), .B1(n13898), .B2(img[631]), .O(
        n16134) );
  AOI22S U18990 ( .A1(n17382), .A2(img[1527]), .B1(n18751), .B2(img[1399]), 
        .O(n16141) );
  AOI22S U18991 ( .A1(n18819), .A2(img[2039]), .B1(n17383), .B2(img[1911]), 
        .O(n16140) );
  INV1S U18992 ( .I(n13789), .O(n18975) );
  AOI22S U18993 ( .A1(n18975), .A2(img[1271]), .B1(n18922), .B2(img[1143]), 
        .O(n16139) );
  AOI22S U18994 ( .A1(n13786), .A2(img[1783]), .B1(n17561), .B2(img[1655]), 
        .O(n16138) );
  AN4S U18995 ( .I1(n16141), .I2(n16140), .I3(n16139), .I4(n16138), .O(n16142)
         );
  ND2S U18996 ( .I1(n16143), .I2(n16142), .O(n20259) );
  AOI22S U18997 ( .A1(n20612), .A2(n13804), .B1(n13846), .B2(n20259), .O(
        n16165) );
  AOI22S U18998 ( .A1(n20102), .A2(img[479]), .B1(n13855), .B2(img[351]), .O(
        n16147) );
  AOI22S U18999 ( .A1(n13788), .A2(img[991]), .B1(n13892), .B2(img[863]), .O(
        n16146) );
  AOI22S U19000 ( .A1(n17197), .A2(img[223]), .B1(n17376), .B2(img[95]), .O(
        n16145) );
  AOI22S U19001 ( .A1(n16348), .A2(img[735]), .B1(n13898), .B2(img[607]), .O(
        n16144) );
  AN4S U19002 ( .I1(n16147), .I2(n16146), .I3(n16145), .I4(n16144), .O(n16153)
         );
  AOI22S U19003 ( .A1(n19193), .A2(img[1503]), .B1(n17827), .B2(img[1375]), 
        .O(n16151) );
  AOI22S U19004 ( .A1(n13841), .A2(img[2015]), .B1(n17383), .B2(img[1887]), 
        .O(n16150) );
  AOI22S U19005 ( .A1(n13853), .A2(img[1247]), .B1(n18974), .B2(img[1119]), 
        .O(n16149) );
  AOI22S U19006 ( .A1(n13867), .A2(img[1759]), .B1(n17550), .B2(img[1631]), 
        .O(n16148) );
  AN4S U19007 ( .I1(n16151), .I2(n16150), .I3(n16149), .I4(n16148), .O(n16152)
         );
  ND2 U19008 ( .I1(n16153), .I2(n16152), .O(n20630) );
  AOI22S U19009 ( .A1(n18681), .A2(img[471]), .B1(n13855), .B2(img[343]), .O(
        n16157) );
  AOI22S U19010 ( .A1(n19649), .A2(img[983]), .B1(n13890), .B2(img[855]), .O(
        n16156) );
  BUF1 U19011 ( .I(n13800), .O(n17218) );
  AOI22S U19012 ( .A1(n17218), .A2(img[215]), .B1(n17376), .B2(img[87]), .O(
        n16155) );
  AOI22S U19013 ( .A1(n16348), .A2(img[727]), .B1(n13797), .B2(img[599]), .O(
        n16154) );
  AN4S U19014 ( .I1(n16157), .I2(n16156), .I3(n16155), .I4(n16154), .O(n16163)
         );
  AOI22S U19015 ( .A1(n19193), .A2(img[1495]), .B1(n18751), .B2(img[1367]), 
        .O(n16161) );
  AOI22S U19016 ( .A1(n17816), .A2(img[2007]), .B1(n17383), .B2(img[1879]), 
        .O(n16160) );
  AOI22S U19017 ( .A1(n16635), .A2(img[1239]), .B1(n18548), .B2(img[1111]), 
        .O(n16159) );
  AOI22S U19018 ( .A1(n13786), .A2(img[1751]), .B1(n17550), .B2(img[1623]), 
        .O(n16158) );
  AN4S U19019 ( .I1(n16161), .I2(n16160), .I3(n16159), .I4(n16158), .O(n16162)
         );
  ND2 U19020 ( .I1(n16163), .I2(n16162), .O(n20607) );
  AOI22S U19021 ( .A1(n20630), .A2(n19914), .B1(n13791), .B2(n20607), .O(
        n16164) );
  AN4S U19022 ( .I1(n16167), .I2(n16166), .I3(n16165), .I4(n16164), .O(n16212)
         );
  ND2 U19023 ( .I1(n16168), .I2(n16212), .O(n16226) );
  INV1S U19024 ( .I(n23973), .O(n16170) );
  NR2 U19025 ( .I1(n23900), .I2(img_size[3]), .O(n16169) );
  BUF1S U19026 ( .I(i_row[3]), .O(n23828) );
  XNR2HS U19027 ( .I1(n23900), .I2(n24332), .O(n23869) );
  INV1S U19028 ( .I(n23869), .O(n23791) );
  XNR2HS U19029 ( .I1(i_row[2]), .I2(n23869), .O(n16176) );
  XOR2HS U19030 ( .I1(i_row[1]), .I2(n23740), .O(n16174) );
  XOR2HS U19031 ( .I1(i_row[0]), .I2(n28555), .O(n16173) );
  ND2S U19032 ( .I1(n16174), .I2(n16173), .O(n16175) );
  XNR2HS U19033 ( .I1(i_col[3]), .I2(n23867), .O(n16179) );
  XNR2HS U19034 ( .I1(i_col[2]), .I2(n23869), .O(n16183) );
  XOR2HS U19035 ( .I1(i_col[1]), .I2(n23740), .O(n16181) );
  XOR2HS U19036 ( .I1(i_col[0]), .I2(n28555), .O(n16180) );
  ND2S U19037 ( .I1(n16181), .I2(n16180), .O(n16182) );
  NR2 U19038 ( .I1(n16183), .I2(n16182), .O(n16184) );
  ND2P U19039 ( .I1(n23601), .I2(n13844), .O(n19700) );
  INV3 U19040 ( .I(n19542), .O(n20371) );
  OR2P U19041 ( .I1(n20969), .I2(n23601), .O(n18132) );
  NR2 U19042 ( .I1(n18141), .I2(n18132), .O(n16187) );
  BUF3 U19043 ( .I(n16187), .O(n19533) );
  AOI22S U19044 ( .A1(n16226), .A2(n20371), .B1(n19533), .B2(n16226), .O(
        n16214) );
  NR2P U19045 ( .I1(n18132), .I2(n18133), .O(n16188) );
  INV2 U19046 ( .I(n22928), .O(n18141) );
  ND2P U19047 ( .I1(n13910), .I2(n18141), .O(n19473) );
  AOI22S U19048 ( .A1(n18681), .A2(img[511]), .B1(n13896), .B2(img[383]), .O(
        n16193) );
  AOI22S U19049 ( .A1(n16515), .A2(img[1023]), .B1(n16048), .B2(img[895]), .O(
        n16192) );
  AOI22S U19050 ( .A1(n17880), .A2(img[255]), .B1(n19642), .B2(img[127]), .O(
        n16191) );
  AOI22S U19051 ( .A1(n13886), .A2(img[767]), .B1(n13797), .B2(img[639]), .O(
        n16190) );
  AN4S U19052 ( .I1(n16193), .I2(n16192), .I3(n16191), .I4(n16190), .O(n16199)
         );
  AOI22S U19053 ( .A1(n19193), .A2(img[1535]), .B1(n18751), .B2(img[1407]), 
        .O(n16197) );
  AOI22S U19054 ( .A1(n19290), .A2(img[2047]), .B1(n22928), .B2(img[1919]), 
        .O(n16196) );
  AOI22S U19055 ( .A1(n17323), .A2(img[1279]), .B1(n18922), .B2(img[1151]), 
        .O(n16195) );
  AOI22S U19056 ( .A1(n13867), .A2(img[1791]), .B1(n17561), .B2(img[1663]), 
        .O(n16194) );
  AN4S U19057 ( .I1(n16197), .I2(n16196), .I3(n16195), .I4(n16194), .O(n16198)
         );
  NR2 U19058 ( .I1(n18141), .I2(n13844), .O(n16200) );
  AOI22S U19059 ( .A1(n19603), .A2(n21259), .B1(n20608), .B2(n22923), .O(
        n16202) );
  ND2S U19060 ( .I1(n20611), .I2(n13839), .O(n16205) );
  ND2S U19061 ( .I1(n20610), .I2(n17875), .O(n16204) );
  ND2S U19062 ( .I1(n16208), .I2(n16207), .O(n16209) );
  NR2 U19063 ( .I1(n16210), .I2(n16209), .O(n16211) );
  INV1S U19064 ( .I(n19608), .O(n17636) );
  AO12 U19065 ( .B1(n16212), .B2(n16211), .A1(n17636), .O(n16215) );
  INV1S U19066 ( .I(n21467), .O(n20383) );
  OR2 U19067 ( .I1(n13822), .I2(n16215), .O(n16263) );
  INV3 U19068 ( .I(n19542), .O(n20314) );
  AN2T U19069 ( .I1(n20314), .I2(n20809), .O(n20223) );
  AOI22S U19070 ( .A1(n20609), .A2(n13839), .B1(n17875), .B2(n20626), .O(
        n16219) );
  AOI22S U19071 ( .A1(n20630), .A2(n19483), .B1(n20187), .B2(n20610), .O(
        n16218) );
  AOI22S U19072 ( .A1(n20612), .A2(n20613), .B1(n17762), .B2(n20624), .O(
        n16217) );
  AOI22S U19073 ( .A1(n20627), .A2(n13830), .B1(n17928), .B2(n20619), .O(
        n16216) );
  AN4S U19074 ( .I1(n16219), .I2(n16218), .I3(n16217), .I4(n16216), .O(n16225)
         );
  AOI22S U19075 ( .A1(n20606), .A2(n20263), .B1(n13847), .B2(n20608), .O(
        n16223) );
  BUF1 U19076 ( .I(n18040), .O(n21061) );
  ND2S U19077 ( .I1(n20628), .I2(n21061), .O(n16222) );
  AOI22S U19078 ( .A1(n20611), .A2(n13846), .B1(n20438), .B2(n20621), .O(
        n16221) );
  AOI22S U19079 ( .A1(n20614), .A2(n13791), .B1(n19914), .B2(n20607), .O(
        n16220) );
  AN4S U19080 ( .I1(n16223), .I2(n16222), .I3(n16221), .I4(n16220), .O(n16224)
         );
  AOI22S U19081 ( .A1(n16226), .A2(n20223), .B1(n16188), .B2(n16260), .O(
        n16262) );
  NR2T U19082 ( .I1(n21237), .I2(n21654), .O(n16255) );
  MOAI1S U19083 ( .A1(n16228), .A2(n15142), .B1(n16227), .B2(n17931), .O(
        n16232) );
  MOAI1S U19084 ( .A1(n16230), .A2(n13945), .B1(n16229), .B2(n21062), .O(
        n16231) );
  NR2 U19085 ( .I1(n16232), .I2(n16231), .O(n16254) );
  INV1S U19086 ( .I(n16233), .O(n16235) );
  AOI22S U19087 ( .A1(n16235), .A2(n20613), .B1(n13791), .B2(n16234), .O(
        n16253) );
  AOI22S U19088 ( .A1(n16237), .A2(n17928), .B1(n16236), .B2(n20969), .O(
        n16252) );
  MOAI1S U19089 ( .A1(n16239), .A2(n13766), .B1(n16238), .B2(n20263), .O(
        n16243) );
  MOAI1S U19090 ( .A1(n16241), .A2(n17656), .B1(n16240), .B2(n18040), .O(
        n16242) );
  NR2 U19091 ( .I1(n16243), .I2(n16242), .O(n16250) );
  AOI22S U19092 ( .A1(n16245), .A2(n13847), .B1(n17875), .B2(n16244), .O(
        n16249) );
  AOI22S U19093 ( .A1(n16247), .A2(n13839), .B1(n13846), .B2(n16246), .O(
        n16248) );
  ND3S U19094 ( .I1(n16250), .I2(n16249), .I3(n16248), .O(n16251) );
  AN4B1S U19095 ( .I1(n16254), .I2(n16253), .I3(n16252), .B1(n16251), .O(
        n20291) );
  AN2 U19096 ( .I1(n21654), .I2(n20291), .O(n20691) );
  ND2S U19097 ( .I1(n21669), .I2(n19603), .O(n16257) );
  ND3HT U19098 ( .I1(n16263), .I2(n16262), .I3(n16261), .O(n22053) );
  AOI22S U19099 ( .A1(n19343), .A2(img[494]), .B1(n13879), .B2(img[366]), .O(
        n16267) );
  AOI22S U19100 ( .A1(n18946), .A2(img[1006]), .B1(n13890), .B2(img[878]), .O(
        n16266) );
  AOI22S U19101 ( .A1(n17377), .A2(img[238]), .B1(n17611), .B2(img[110]), .O(
        n16265) );
  BUF1 U19102 ( .I(n15568), .O(n17835) );
  AOI22S U19103 ( .A1(n17835), .A2(img[750]), .B1(n13837), .B2(img[622]), .O(
        n16264) );
  AN4S U19104 ( .I1(n16267), .I2(n16266), .I3(n16265), .I4(n16264), .O(n16273)
         );
  AOI22S U19105 ( .A1(n15630), .A2(img[1518]), .B1(n17862), .B2(img[1390]), 
        .O(n16271) );
  BUF6CK U19106 ( .I(n15080), .O(n17863) );
  AOI22S U19107 ( .A1(n17886), .A2(img[2030]), .B1(n17863), .B2(img[1902]), 
        .O(n16270) );
  AOI22S U19108 ( .A1(n17347), .A2(img[1262]), .B1(n17840), .B2(img[1134]), 
        .O(n16269) );
  AOI22S U19109 ( .A1(n19023), .A2(img[1774]), .B1(n17561), .B2(img[1646]), 
        .O(n16268) );
  AN4S U19110 ( .I1(n16271), .I2(n16270), .I3(n16269), .I4(n16268), .O(n16272)
         );
  AOI22S U19111 ( .A1(n19343), .A2(img[430]), .B1(n13855), .B2(img[302]), .O(
        n16278) );
  AOI22S U19112 ( .A1(n18935), .A2(img[942]), .B1(n15653), .B2(img[814]), .O(
        n16277) );
  AOI22S U19113 ( .A1(n18796), .A2(img[174]), .B1(n17611), .B2(img[46]), .O(
        n16276) );
  AOI22S U19114 ( .A1(n13875), .A2(img[686]), .B1(n13837), .B2(img[558]), .O(
        n16275) );
  AOI22S U19115 ( .A1(n19193), .A2(img[1454]), .B1(n13798), .B2(img[1326]), 
        .O(n16282) );
  AOI22S U19116 ( .A1(n18958), .A2(img[1966]), .B1(n17863), .B2(img[1838]), 
        .O(n16281) );
  AOI22S U19117 ( .A1(n18923), .A2(img[1198]), .B1(n17712), .B2(img[1070]), 
        .O(n16280) );
  AOI22S U19118 ( .A1(n19023), .A2(img[1710]), .B1(n13832), .B2(img[1582]), 
        .O(n16279) );
  ND2P U19119 ( .I1(n16284), .I2(n16283), .O(n20592) );
  AOI22S U19120 ( .A1(n20593), .A2(n13839), .B1(n17875), .B2(n20592), .O(
        n16347) );
  AOI22S U19121 ( .A1(n13825), .A2(img[438]), .B1(n13859), .B2(img[310]), .O(
        n16288) );
  AOI22S U19122 ( .A1(n19037), .A2(img[950]), .B1(n13890), .B2(img[822]), .O(
        n16287) );
  AOI22S U19123 ( .A1(n19266), .A2(img[182]), .B1(n17611), .B2(img[54]), .O(
        n16286) );
  AOI22S U19124 ( .A1(n13875), .A2(img[694]), .B1(n13797), .B2(img[566]), .O(
        n16285) );
  AN4S U19125 ( .I1(n16288), .I2(n16287), .I3(n16286), .I4(n16285), .O(n16295)
         );
  AOI22S U19126 ( .A1(n13823), .A2(img[1462]), .B1(n16127), .B2(img[1334]), 
        .O(n16293) );
  AOI22S U19127 ( .A1(n13841), .A2(img[1974]), .B1(n17863), .B2(img[1846]), 
        .O(n16292) );
  AOI22S U19128 ( .A1(n17347), .A2(img[1206]), .B1(n13802), .B2(img[1078]), 
        .O(n16291) );
  AOI22S U19129 ( .A1(n19215), .A2(img[1718]), .B1(n13796), .B2(img[1590]), 
        .O(n16290) );
  AN4S U19130 ( .I1(n16293), .I2(n16292), .I3(n16291), .I4(n16290), .O(n16294)
         );
  ND2P U19131 ( .I1(n16295), .I2(n16294), .O(n20569) );
  AOI22S U19132 ( .A1(n19343), .A2(img[486]), .B1(n19709), .B2(img[358]), .O(
        n16299) );
  AOI22S U19133 ( .A1(n14822), .A2(img[998]), .B1(n16048), .B2(img[870]), .O(
        n16298) );
  BUF1 U19134 ( .I(n13800), .O(n17729) );
  AOI22S U19135 ( .A1(n17729), .A2(img[230]), .B1(n17611), .B2(img[102]), .O(
        n16297) );
  AOI22S U19136 ( .A1(n17730), .A2(img[742]), .B1(n13898), .B2(img[614]), .O(
        n16296) );
  AN4S U19137 ( .I1(n16299), .I2(n16298), .I3(n16297), .I4(n16296), .O(n16305)
         );
  AOI22S U19138 ( .A1(n19193), .A2(img[1510]), .B1(n17862), .B2(img[1382]), 
        .O(n16303) );
  AOI22S U19139 ( .A1(n13803), .A2(img[2022]), .B1(n17863), .B2(img[1894]), 
        .O(n16302) );
  AOI22S U19140 ( .A1(n16799), .A2(img[1254]), .B1(n13802), .B2(img[1126]), 
        .O(n16301) );
  AOI22S U19141 ( .A1(n13786), .A2(img[1766]), .B1(n17561), .B2(img[1638]), 
        .O(n16300) );
  AN4S U19142 ( .I1(n16303), .I2(n16302), .I3(n16301), .I4(n16300), .O(n16304)
         );
  ND2 U19143 ( .I1(n16305), .I2(n16304), .O(n20588) );
  AOI22S U19144 ( .A1(n20569), .A2(n20187), .B1(n21062), .B2(n20588), .O(
        n16443) );
  AOI22S U19145 ( .A1(n19343), .A2(img[422]), .B1(n19709), .B2(img[294]), .O(
        n16309) );
  AOI22S U19146 ( .A1(n16515), .A2(img[934]), .B1(n13893), .B2(img[806]), .O(
        n16308) );
  AOI22S U19147 ( .A1(n17377), .A2(img[166]), .B1(n17611), .B2(img[38]), .O(
        n16307) );
  AOI22S U19148 ( .A1(n19641), .A2(img[678]), .B1(n13797), .B2(img[550]), .O(
        n16306) );
  AN4S U19149 ( .I1(n16309), .I2(n16308), .I3(n16307), .I4(n16306), .O(n16315)
         );
  AOI22S U19150 ( .A1(n19193), .A2(img[1446]), .B1(n17827), .B2(img[1318]), 
        .O(n16313) );
  AOI22S U19151 ( .A1(n20104), .A2(img[1958]), .B1(n17863), .B2(img[1830]), 
        .O(n16312) );
  AOI22S U19152 ( .A1(n14392), .A2(img[1190]), .B1(n17745), .B2(img[1062]), 
        .O(n16311) );
  AOI22S U19153 ( .A1(n19215), .A2(img[1702]), .B1(n17561), .B2(img[1574]), 
        .O(n16310) );
  AN4S U19154 ( .I1(n16313), .I2(n16312), .I3(n16311), .I4(n16310), .O(n16314)
         );
  ND2 U19155 ( .I1(n16315), .I2(n16314), .O(n20577) );
  AOI22S U19156 ( .A1(n19343), .A2(img[406]), .B1(n13896), .B2(img[278]), .O(
        n16319) );
  AOI22S U19157 ( .A1(n18148), .A2(img[918]), .B1(n13892), .B2(img[790]), .O(
        n16318) );
  AOI22S U19158 ( .A1(n17218), .A2(img[150]), .B1(n17611), .B2(img[22]), .O(
        n16317) );
  AOI22S U19159 ( .A1(n13784), .A2(img[662]), .B1(n13898), .B2(img[534]), .O(
        n16316) );
  AN4S U19160 ( .I1(n16319), .I2(n16318), .I3(n16317), .I4(n16316), .O(n16325)
         );
  AOI22S U19161 ( .A1(n19193), .A2(img[1430]), .B1(n17827), .B2(img[1302]), 
        .O(n16323) );
  AOI22S U19162 ( .A1(n13803), .A2(img[1942]), .B1(n17863), .B2(img[1814]), 
        .O(n16322) );
  AOI22S U19163 ( .A1(n13853), .A2(img[1174]), .B1(n18922), .B2(img[1046]), 
        .O(n16321) );
  AOI22S U19164 ( .A1(n13786), .A2(img[1686]), .B1(n17561), .B2(img[1558]), 
        .O(n16320) );
  AN4S U19165 ( .I1(n16323), .I2(n16322), .I3(n16321), .I4(n16320), .O(n16324)
         );
  AOI22S U19166 ( .A1(n20577), .A2(n20613), .B1(n17762), .B2(n20570), .O(
        n16445) );
  AOI22S U19167 ( .A1(n15506), .A2(img[398]), .B1(n15691), .B2(img[270]), .O(
        n16330) );
  AOI22S U19168 ( .A1(n16515), .A2(img[910]), .B1(n13861), .B2(img[782]), .O(
        n16329) );
  AOI22S U19169 ( .A1(n13800), .A2(img[142]), .B1(n17376), .B2(img[14]), .O(
        n16328) );
  AOI22S U19170 ( .A1(n19252), .A2(img[654]), .B1(n13797), .B2(img[526]), .O(
        n16327) );
  AN4S U19171 ( .I1(n16330), .I2(n16329), .I3(n16328), .I4(n16327), .O(n16336)
         );
  AOI22S U19172 ( .A1(n19193), .A2(img[1422]), .B1(n13798), .B2(img[1294]), 
        .O(n16334) );
  AOI22S U19173 ( .A1(n13803), .A2(img[1934]), .B1(n17863), .B2(img[1806]), 
        .O(n16333) );
  AOI22S U19174 ( .A1(n17347), .A2(img[1166]), .B1(n17767), .B2(img[1038]), 
        .O(n16332) );
  AOI22S U19175 ( .A1(n19023), .A2(img[1678]), .B1(n13796), .B2(img[1550]), 
        .O(n16331) );
  AN4S U19176 ( .I1(n16334), .I2(n16333), .I3(n16332), .I4(n16331), .O(n16335)
         );
  AOI22S U19177 ( .A1(n19343), .A2(img[446]), .B1(n13859), .B2(img[318]), .O(
        n16340) );
  AOI22S U19178 ( .A1(n18946), .A2(img[958]), .B1(n13893), .B2(img[830]), .O(
        n16339) );
  BUF1 U19179 ( .I(n13800), .O(n17811) );
  AOI22S U19180 ( .A1(n17811), .A2(img[190]), .B1(n19388), .B2(img[62]), .O(
        n16338) );
  AOI22S U19181 ( .A1(n16348), .A2(img[702]), .B1(n13837), .B2(img[574]), .O(
        n16337) );
  AN4S U19182 ( .I1(n16340), .I2(n16339), .I3(n16338), .I4(n16337), .O(n16346)
         );
  AOI22S U19183 ( .A1(n13823), .A2(img[1470]), .B1(n17862), .B2(img[1342]), 
        .O(n16344) );
  AOI22S U19184 ( .A1(n17816), .A2(img[1982]), .B1(n17863), .B2(img[1854]), 
        .O(n16343) );
  AOI22S U19185 ( .A1(n13783), .A2(img[1214]), .B1(n13787), .B2(img[1086]), 
        .O(n16342) );
  AOI22S U19186 ( .A1(n13870), .A2(img[1726]), .B1(n13794), .B2(img[1598]), 
        .O(n16341) );
  AOI22S U19187 ( .A1(n20573), .A2(n13830), .B1(n17928), .B2(n20579), .O(
        n16444) );
  AN4S U19188 ( .I1(n16347), .I2(n16443), .I3(n16445), .I4(n16444), .O(n16426)
         );
  AOI22S U19189 ( .A1(n13785), .A2(img[462]), .B1(n13855), .B2(img[334]), .O(
        n16352) );
  AOI22S U19190 ( .A1(n18946), .A2(img[974]), .B1(n13893), .B2(img[846]), .O(
        n16351) );
  BUF1 U19191 ( .I(n13800), .O(n17788) );
  AOI22S U19192 ( .A1(n17788), .A2(img[206]), .B1(n17611), .B2(img[78]), .O(
        n16350) );
  AOI22S U19193 ( .A1(n16348), .A2(img[718]), .B1(n13837), .B2(img[590]), .O(
        n16349) );
  AN4S U19194 ( .I1(n16352), .I2(n16351), .I3(n16350), .I4(n16349), .O(n16359)
         );
  AOI22S U19195 ( .A1(n19193), .A2(img[1486]), .B1(n16353), .B2(img[1358]), 
        .O(n16357) );
  AOI22S U19196 ( .A1(n17864), .A2(img[1998]), .B1(n17863), .B2(img[1870]), 
        .O(n16356) );
  AOI22S U19197 ( .A1(n15315), .A2(img[1230]), .B1(n13802), .B2(img[1102]), 
        .O(n16355) );
  AOI22S U19198 ( .A1(n19036), .A2(img[1742]), .B1(n13794), .B2(img[1614]), 
        .O(n16354) );
  AN4S U19199 ( .I1(n16357), .I2(n16356), .I3(n16355), .I4(n16354), .O(n16358)
         );
  AOI22S U19200 ( .A1(n20032), .A2(img[390]), .B1(n13879), .B2(img[262]), .O(
        n16363) );
  AOI22S U19201 ( .A1(n16515), .A2(img[902]), .B1(n15653), .B2(img[774]), .O(
        n16362) );
  AOI22S U19202 ( .A1(n17488), .A2(img[134]), .B1(n19388), .B2(img[6]), .O(
        n16361) );
  AOI22S U19203 ( .A1(n19641), .A2(img[646]), .B1(n13797), .B2(img[518]), .O(
        n16360) );
  AN4S U19204 ( .I1(n16363), .I2(n16362), .I3(n16361), .I4(n16360), .O(n16370)
         );
  AOI22S U19205 ( .A1(n19193), .A2(img[1414]), .B1(n19001), .B2(img[1286]), 
        .O(n16368) );
  AOI22S U19206 ( .A1(n13803), .A2(img[1926]), .B1(n17863), .B2(img[1798]), 
        .O(n16367) );
  AOI22S U19207 ( .A1(n18778), .A2(img[1158]), .B1(n17745), .B2(img[1030]), 
        .O(n16366) );
  AOI22S U19208 ( .A1(n15751), .A2(img[1670]), .B1(n13794), .B2(img[1542]), 
        .O(n16365) );
  AOI22S U19209 ( .A1(n20595), .A2(n20439), .B1(n13847), .B2(n20578), .O(
        n16425) );
  AOI22S U19210 ( .A1(n15506), .A2(img[454]), .B1(n13896), .B2(img[326]), .O(
        n16374) );
  AOI22S U19211 ( .A1(n18148), .A2(img[966]), .B1(n13877), .B2(img[838]), .O(
        n16373) );
  AOI22S U19212 ( .A1(n17811), .A2(img[198]), .B1(n20103), .B2(img[70]), .O(
        n16372) );
  AOI22S U19213 ( .A1(n19252), .A2(img[710]), .B1(n13837), .B2(img[582]), .O(
        n16371) );
  AN4S U19214 ( .I1(n16374), .I2(n16373), .I3(n16372), .I4(n16371), .O(n16381)
         );
  AOI22S U19215 ( .A1(n19193), .A2(img[1478]), .B1(n13798), .B2(img[1350]), 
        .O(n16379) );
  AOI22S U19216 ( .A1(n13801), .A2(img[1990]), .B1(n17863), .B2(img[1862]), 
        .O(n16378) );
  AOI22S U19217 ( .A1(n13853), .A2(img[1222]), .B1(n15800), .B2(img[1094]), 
        .O(n16377) );
  AOI22S U19218 ( .A1(n13786), .A2(img[1734]), .B1(n17561), .B2(img[1606]), 
        .O(n16376) );
  AN4S U19219 ( .I1(n16379), .I2(n16378), .I3(n16377), .I4(n16376), .O(n16380)
         );
  BUF1 U19220 ( .I(n18040), .O(n20580) );
  AOI22S U19221 ( .A1(n13883), .A2(img[414]), .B1(n13896), .B2(img[286]), .O(
        n16385) );
  AOI22S U19222 ( .A1(n18935), .A2(img[926]), .B1(n13893), .B2(img[798]), .O(
        n16384) );
  AOI22S U19223 ( .A1(n19266), .A2(img[158]), .B1(n17611), .B2(img[30]), .O(
        n16383) );
  AOI22S U19224 ( .A1(n19641), .A2(img[670]), .B1(n13837), .B2(img[542]), .O(
        n16382) );
  AN4S U19225 ( .I1(n16385), .I2(n16384), .I3(n16383), .I4(n16382), .O(n16391)
         );
  AOI22S U19226 ( .A1(n19193), .A2(img[1438]), .B1(n13798), .B2(img[1310]), 
        .O(n16389) );
  AOI22S U19227 ( .A1(n18819), .A2(img[1950]), .B1(n17863), .B2(img[1822]), 
        .O(n16388) );
  AOI22S U19228 ( .A1(n13783), .A2(img[1182]), .B1(n17745), .B2(img[1054]), 
        .O(n16387) );
  AOI22S U19229 ( .A1(n16075), .A2(img[1694]), .B1(n13796), .B2(img[1566]), 
        .O(n16386) );
  AN4S U19230 ( .I1(n16389), .I2(n16388), .I3(n16387), .I4(n16386), .O(n16390)
         );
  AOI22S U19231 ( .A1(n18681), .A2(img[502]), .B1(n13879), .B2(img[374]), .O(
        n16395) );
  AOI22S U19232 ( .A1(n13788), .A2(img[1014]), .B1(n13861), .B2(img[886]), .O(
        n16394) );
  AOI22S U19233 ( .A1(n19266), .A2(img[246]), .B1(n17611), .B2(img[118]), .O(
        n16393) );
  AOI22S U19234 ( .A1(n16348), .A2(img[758]), .B1(n13837), .B2(img[630]), .O(
        n16392) );
  AN4S U19235 ( .I1(n16395), .I2(n16394), .I3(n16393), .I4(n16392), .O(n16401)
         );
  AOI22S U19236 ( .A1(n17382), .A2(img[1526]), .B1(n13798), .B2(img[1398]), 
        .O(n16399) );
  AOI22S U19237 ( .A1(n18958), .A2(img[2038]), .B1(n17863), .B2(img[1910]), 
        .O(n16398) );
  AOI22S U19238 ( .A1(n18824), .A2(img[1270]), .B1(n19955), .B2(img[1142]), 
        .O(n16397) );
  AOI22S U19239 ( .A1(n19036), .A2(img[1782]), .B1(n17561), .B2(img[1654]), 
        .O(n16396) );
  AN4S U19240 ( .I1(n16399), .I2(n16398), .I3(n16397), .I4(n16396), .O(n16400)
         );
  AOI22S U19241 ( .A1(n20594), .A2(n13804), .B1(n13846), .B2(n19929), .O(
        n16423) );
  AOI22S U19242 ( .A1(n13785), .A2(img[478]), .B1(n13855), .B2(img[350]), .O(
        n16405) );
  AOI22S U19243 ( .A1(n18988), .A2(img[990]), .B1(n16048), .B2(img[862]), .O(
        n16404) );
  BUF1 U19244 ( .I(n13800), .O(n17857) );
  AOI22S U19245 ( .A1(n17857), .A2(img[222]), .B1(n17611), .B2(img[94]), .O(
        n16403) );
  AOI22S U19246 ( .A1(n19641), .A2(img[734]), .B1(n13837), .B2(img[606]), .O(
        n16402) );
  AN4S U19247 ( .I1(n16405), .I2(n16404), .I3(n16403), .I4(n16402), .O(n16411)
         );
  AOI22S U19248 ( .A1(n13874), .A2(img[1502]), .B1(n16127), .B2(img[1374]), 
        .O(n16409) );
  AOI22S U19249 ( .A1(n17778), .A2(img[2014]), .B1(n17863), .B2(img[1886]), 
        .O(n16408) );
  AOI22S U19250 ( .A1(n18897), .A2(img[1246]), .B1(n17865), .B2(img[1118]), 
        .O(n16407) );
  AOI22S U19251 ( .A1(n19023), .A2(img[1758]), .B1(n13794), .B2(img[1630]), 
        .O(n16406) );
  AN4S U19252 ( .I1(n16409), .I2(n16408), .I3(n16407), .I4(n16406), .O(n16410)
         );
  AOI22S U19253 ( .A1(n13876), .A2(img[470]), .B1(n19709), .B2(img[342]), .O(
        n16415) );
  AOI22S U19254 ( .A1(n18911), .A2(img[982]), .B1(n13893), .B2(img[854]), .O(
        n16414) );
  AOI22S U19255 ( .A1(n17857), .A2(img[214]), .B1(n19388), .B2(img[86]), .O(
        n16413) );
  AOI22S U19256 ( .A1(n19641), .A2(img[726]), .B1(n13797), .B2(img[598]), .O(
        n16412) );
  AN4S U19257 ( .I1(n16415), .I2(n16414), .I3(n16413), .I4(n16412), .O(n16421)
         );
  AOI22S U19258 ( .A1(n20109), .A2(img[1494]), .B1(n17862), .B2(img[1366]), 
        .O(n16419) );
  AOI22S U19259 ( .A1(n19411), .A2(img[2006]), .B1(n17863), .B2(img[1878]), 
        .O(n16418) );
  AOI22S U19260 ( .A1(n17359), .A2(img[1238]), .B1(n17865), .B2(img[1110]), 
        .O(n16417) );
  AOI22S U19261 ( .A1(n19036), .A2(img[1750]), .B1(n13794), .B2(img[1622]), 
        .O(n16416) );
  AN4S U19262 ( .I1(n16419), .I2(n16418), .I3(n16417), .I4(n16416), .O(n16420)
         );
  ND2 U19263 ( .I1(n16421), .I2(n16420), .O(n19930) );
  AOI22S U19264 ( .A1(n20581), .A2(n19914), .B1(n17938), .B2(n19930), .O(
        n16422) );
  AN4 U19265 ( .I1(n16425), .I2(n16424), .I3(n16423), .I4(n16422), .O(n16449)
         );
  ND2S U19266 ( .I1(n16426), .I2(n16449), .O(n16463) );
  AOI22S U19267 ( .A1(n16463), .A2(n20371), .B1(n19533), .B2(n16463), .O(
        n16451) );
  AOI22S U19268 ( .A1(n13825), .A2(img[510]), .B1(n13858), .B2(img[382]), .O(
        n16430) );
  AOI22S U19269 ( .A1(n17880), .A2(img[254]), .B1(n19642), .B2(img[126]), .O(
        n16429) );
  AOI22S U19270 ( .A1(n18988), .A2(img[1022]), .B1(n13890), .B2(img[894]), .O(
        n16428) );
  AOI22S U19271 ( .A1(n13886), .A2(img[766]), .B1(n13898), .B2(img[638]), .O(
        n16427) );
  AN4S U19272 ( .I1(n16430), .I2(n16429), .I3(n16428), .I4(n16427), .O(n16437)
         );
  AOI22S U19273 ( .A1(n13783), .A2(img[1278]), .B1(n17885), .B2(img[1150]), 
        .O(n16435) );
  AOI22S U19274 ( .A1(n15809), .A2(img[1790]), .B1(n17561), .B2(img[1662]), 
        .O(n16434) );
  AOI22S U19275 ( .A1(n13823), .A2(img[1534]), .B1(n19182), .B2(img[1406]), 
        .O(n16433) );
  AOI22S U19276 ( .A1(n13801), .A2(img[2046]), .B1(n22928), .B2(img[1918]), 
        .O(n16432) );
  AN4S U19277 ( .I1(n16435), .I2(n16434), .I3(n16433), .I4(n16432), .O(n16436)
         );
  ND2 U19278 ( .I1(n16437), .I2(n16436), .O(n19939) );
  AOI22S U19279 ( .A1(n19603), .A2(n21254), .B1(n19939), .B2(n22923), .O(
        n16439) );
  ND2S U19280 ( .I1(n16439), .I2(n16438), .O(n16440) );
  AOI12HS U19281 ( .B1(n16463), .B2(n20364), .A1(n16440), .O(n16450) );
  ND2S U19282 ( .I1(n20593), .I2(n13839), .O(n16442) );
  ND2S U19283 ( .I1(n20592), .I2(n17875), .O(n16441) );
  ND3S U19284 ( .I1(n16443), .I2(n16442), .I3(n16441), .O(n16447) );
  ND2S U19285 ( .I1(n16445), .I2(n16444), .O(n16446) );
  NR2 U19286 ( .I1(n16447), .I2(n16446), .O(n16448) );
  AO12 U19287 ( .B1(n16449), .B2(n16448), .A1(n17636), .O(n16452) );
  ND2T U19288 ( .I1(n21804), .I2(n20809), .O(n29503) );
  AOI22S U19289 ( .A1(n20588), .A2(n13839), .B1(n17875), .B2(n20577), .O(
        n16456) );
  AOI22S U19290 ( .A1(n20581), .A2(n19483), .B1(n20187), .B2(n20592), .O(
        n16455) );
  AOI22S U19291 ( .A1(n20594), .A2(n20613), .B1(n17762), .B2(n20573), .O(
        n16454) );
  AOI22S U19292 ( .A1(n20578), .A2(n13830), .B1(n17928), .B2(n20569), .O(
        n16453) );
  AN4S U19293 ( .I1(n16456), .I2(n16455), .I3(n16454), .I4(n16453), .O(n16462)
         );
  AOI22S U19294 ( .A1(n20585), .A2(n20439), .B1(n13847), .B2(n19939), .O(
        n16460) );
  ND2S U19295 ( .I1(n20579), .I2(n20629), .O(n16459) );
  AOI22S U19296 ( .A1(n20593), .A2(n13846), .B1(n20438), .B2(n20570), .O(
        n16458) );
  AOI22S U19297 ( .A1(n20595), .A2(n13791), .B1(n13835), .B2(n19930), .O(
        n16457) );
  AN4S U19298 ( .I1(n16460), .I2(n16459), .I3(n16458), .I4(n16457), .O(n16461)
         );
  ND2S U19299 ( .I1(n16462), .I2(n16461), .O(n16502) );
  AOI22S U19300 ( .A1(n16463), .A2(n20223), .B1(n16188), .B2(n16502), .O(
        n16504) );
  AOI22S U19301 ( .A1(n19818), .A2(n19929), .B1(n19929), .B2(n22923), .O(
        n16500) );
  INV1S U19302 ( .I(n19700), .O(n16464) );
  AN2 U19303 ( .I1(n19603), .I2(n21654), .O(n17686) );
  INV1S U19304 ( .I(n16465), .O(n16469) );
  INV1S U19305 ( .I(n16466), .O(n16467) );
  MOAI1 U19306 ( .A1(n16469), .A2(n16468), .B1(n16467), .B2(n13830), .O(n16473) );
  MOAI1S U19307 ( .A1(n16471), .A2(n13766), .B1(n16470), .B2(n13839), .O(
        n16472) );
  NR2 U19308 ( .I1(n16473), .I2(n16472), .O(n16480) );
  AOI22S U19309 ( .A1(n16475), .A2(n19914), .B1(n17928), .B2(n16474), .O(
        n16479) );
  AOI22S U19310 ( .A1(n16477), .A2(n13846), .B1(n13791), .B2(n16476), .O(
        n16478) );
  MOAI1S U19311 ( .A1(n16482), .A2(n17656), .B1(n16481), .B2(n20969), .O(
        n16487) );
  INV1S U19312 ( .I(n16483), .O(n16484) );
  INV1S U19313 ( .I(n16488), .O(n16489) );
  AOI22S U19314 ( .A1(n16490), .A2(n20263), .B1(n13847), .B2(n16489), .O(
        n16495) );
  INV1S U19315 ( .I(n16491), .O(n16492) );
  AOI22S U19316 ( .A1(n16493), .A2(n19483), .B1(n20963), .B2(n16492), .O(
        n16494) );
  AOI22S U19317 ( .A1(n20252), .A2(n21254), .B1(n17686), .B2(n20685), .O(
        n16499) );
  ND2S U19318 ( .I1(n16500), .I2(n16499), .O(n16501) );
  AOI12HS U19319 ( .B1(n16502), .B2(n19533), .A1(n16501), .O(n16503) );
  AOI22S U19320 ( .A1(n20102), .A2(img[493]), .B1(n13855), .B2(img[365]), .O(
        n16508) );
  AOI22S U19321 ( .A1(n14505), .A2(img[1005]), .B1(n13880), .B2(img[877]), .O(
        n16507) );
  AOI22S U19322 ( .A1(n17377), .A2(img[237]), .B1(n17376), .B2(img[109]), .O(
        n16506) );
  AOI22S U19323 ( .A1(n19641), .A2(img[749]), .B1(n13797), .B2(img[621]), .O(
        n16505) );
  AOI22S U19324 ( .A1(n17382), .A2(img[1517]), .B1(n19182), .B2(img[1389]), 
        .O(n16512) );
  AOI22S U19325 ( .A1(n17515), .A2(img[2029]), .B1(n17383), .B2(img[1901]), 
        .O(n16511) );
  AOI22S U19326 ( .A1(n17323), .A2(img[1261]), .B1(n17767), .B2(img[1133]), 
        .O(n16510) );
  AOI22S U19327 ( .A1(n18885), .A2(img[1773]), .B1(n18201), .B2(img[1645]), 
        .O(n16509) );
  AN4S U19328 ( .I1(n16512), .I2(n16511), .I3(n16510), .I4(n16509), .O(n16513)
         );
  AOI22S U19329 ( .A1(n19343), .A2(img[429]), .B1(n13858), .B2(img[301]), .O(
        n16520) );
  AOI22S U19330 ( .A1(n17810), .A2(img[941]), .B1(n16048), .B2(img[813]), .O(
        n16519) );
  AOI22S U19331 ( .A1(n17271), .A2(img[173]), .B1(n17376), .B2(img[45]), .O(
        n16518) );
  AOI22S U19332 ( .A1(n19326), .A2(img[685]), .B1(n13797), .B2(img[557]), .O(
        n16517) );
  AN4S U19333 ( .I1(n16520), .I2(n16519), .I3(n16518), .I4(n16517), .O(n16526)
         );
  AOI22S U19334 ( .A1(n20109), .A2(img[1453]), .B1(n13845), .B2(img[1325]), 
        .O(n16524) );
  AOI22S U19335 ( .A1(n18773), .A2(img[1965]), .B1(n17383), .B2(img[1837]), 
        .O(n16523) );
  INV1S U19336 ( .I(n13789), .O(n17312) );
  AOI22S U19337 ( .A1(n17312), .A2(img[1197]), .B1(n17276), .B2(img[1069]), 
        .O(n16522) );
  AOI22S U19338 ( .A1(n13786), .A2(img[1709]), .B1(n19416), .B2(img[1581]), 
        .O(n16521) );
  AN4S U19339 ( .I1(n16524), .I2(n16523), .I3(n16522), .I4(n16521), .O(n16525)
         );
  ND2P U19340 ( .I1(n16526), .I2(n16525), .O(n20543) );
  AOI22S U19341 ( .A1(n20544), .A2(n13839), .B1(n17875), .B2(n20543), .O(
        n16590) );
  AOI22S U19342 ( .A1(n20032), .A2(img[437]), .B1(n13858), .B2(img[309]), .O(
        n16530) );
  AOI22S U19343 ( .A1(n18946), .A2(img[949]), .B1(n13889), .B2(img[821]), .O(
        n16529) );
  AOI22S U19344 ( .A1(n17534), .A2(img[181]), .B1(n17376), .B2(img[53]), .O(
        n16528) );
  AOI22S U19345 ( .A1(n13875), .A2(img[693]), .B1(n13797), .B2(img[565]), .O(
        n16527) );
  AOI22S U19346 ( .A1(n17382), .A2(img[1461]), .B1(n19182), .B2(img[1333]), 
        .O(n16534) );
  AOI22S U19347 ( .A1(n13833), .A2(img[1973]), .B1(n17383), .B2(img[1845]), 
        .O(n16533) );
  AOI22S U19348 ( .A1(n16635), .A2(img[1205]), .B1(n19647), .B2(img[1077]), 
        .O(n16532) );
  AOI22S U19349 ( .A1(n19023), .A2(img[1717]), .B1(n18201), .B2(img[1589]), 
        .O(n16531) );
  AN4S U19350 ( .I1(n16534), .I2(n16533), .I3(n16532), .I4(n16531), .O(n16535)
         );
  AOI22S U19351 ( .A1(n18681), .A2(img[485]), .B1(n13855), .B2(img[357]), .O(
        n16540) );
  AOI22S U19352 ( .A1(n18946), .A2(img[997]), .B1(n13893), .B2(img[869]), .O(
        n16539) );
  AOI22S U19353 ( .A1(n17197), .A2(img[229]), .B1(n17376), .B2(img[101]), .O(
        n16538) );
  AOI22S U19354 ( .A1(n17730), .A2(img[741]), .B1(n13837), .B2(img[613]), .O(
        n16537) );
  AOI22S U19355 ( .A1(n17382), .A2(img[1509]), .B1(n13798), .B2(img[1381]), 
        .O(n16544) );
  AOI22S U19356 ( .A1(n13801), .A2(img[2021]), .B1(n17383), .B2(img[1893]), 
        .O(n16543) );
  AOI22S U19357 ( .A1(n15315), .A2(img[1253]), .B1(n17840), .B2(img[1125]), 
        .O(n16542) );
  AOI22S U19358 ( .A1(n19036), .A2(img[1765]), .B1(n18201), .B2(img[1637]), 
        .O(n16541) );
  AN4S U19359 ( .I1(n16544), .I2(n16543), .I3(n16542), .I4(n16541), .O(n16545)
         );
  AOI22S U19360 ( .A1(n20551), .A2(n20963), .B1(n21062), .B2(n20542), .O(
        n16589) );
  AOI22S U19361 ( .A1(n13825), .A2(img[421]), .B1(n13858), .B2(img[293]), .O(
        n16550) );
  AOI22S U19362 ( .A1(n14505), .A2(img[933]), .B1(n13893), .B2(img[805]), .O(
        n16549) );
  AOI22S U19363 ( .A1(n19289), .A2(img[165]), .B1(n17376), .B2(img[37]), .O(
        n16548) );
  AOI22S U19364 ( .A1(n13875), .A2(img[677]), .B1(n13837), .B2(img[549]), .O(
        n16547) );
  AN4S U19365 ( .I1(n16550), .I2(n16549), .I3(n16548), .I4(n16547), .O(n16556)
         );
  AOI22S U19366 ( .A1(n19193), .A2(img[1445]), .B1(n13845), .B2(img[1317]), 
        .O(n16554) );
  AOI22S U19367 ( .A1(n17793), .A2(img[1957]), .B1(n17383), .B2(img[1829]), 
        .O(n16553) );
  AOI22S U19368 ( .A1(n17336), .A2(img[1189]), .B1(n13787), .B2(img[1061]), 
        .O(n16552) );
  AOI22S U19369 ( .A1(n15809), .A2(img[1701]), .B1(n13794), .B2(img[1573]), 
        .O(n16551) );
  AN4S U19370 ( .I1(n16554), .I2(n16553), .I3(n16552), .I4(n16551), .O(n16555)
         );
  AOI22S U19371 ( .A1(n13825), .A2(img[405]), .B1(n13858), .B2(img[277]), .O(
        n16560) );
  AOI22S U19372 ( .A1(n17810), .A2(img[917]), .B1(n13877), .B2(img[789]), .O(
        n16559) );
  AOI22S U19373 ( .A1(n17330), .A2(img[149]), .B1(n17376), .B2(img[21]), .O(
        n16558) );
  AOI22S U19374 ( .A1(n16348), .A2(img[661]), .B1(n13797), .B2(img[533]), .O(
        n16557) );
  AN4S U19375 ( .I1(n16560), .I2(n16559), .I3(n16558), .I4(n16557), .O(n16566)
         );
  AOI22S U19376 ( .A1(n19193), .A2(img[1429]), .B1(n17862), .B2(img[1301]), 
        .O(n16564) );
  AOI22S U19377 ( .A1(n20104), .A2(img[1941]), .B1(n17383), .B2(img[1813]), 
        .O(n16563) );
  AOI22S U19378 ( .A1(n17336), .A2(img[1173]), .B1(n18922), .B2(img[1045]), 
        .O(n16562) );
  AOI22S U19379 ( .A1(n19215), .A2(img[1685]), .B1(n17550), .B2(img[1557]), 
        .O(n16561) );
  AN4S U19380 ( .I1(n16564), .I2(n16563), .I3(n16562), .I4(n16561), .O(n16565)
         );
  AOI22S U19381 ( .A1(n20557), .A2(n20613), .B1(n17762), .B2(n20552), .O(
        n16588) );
  AOI22S U19382 ( .A1(n13883), .A2(img[397]), .B1(n13858), .B2(img[269]), .O(
        n16570) );
  AOI22S U19383 ( .A1(n18946), .A2(img[909]), .B1(n13893), .B2(img[781]), .O(
        n16569) );
  AOI22S U19384 ( .A1(n17249), .A2(img[141]), .B1(n17376), .B2(img[13]), .O(
        n16568) );
  AOI22S U19385 ( .A1(n13875), .A2(img[653]), .B1(n13797), .B2(img[525]), .O(
        n16567) );
  AOI22S U19386 ( .A1(n19193), .A2(img[1421]), .B1(n17862), .B2(img[1293]), 
        .O(n16574) );
  AOI22S U19387 ( .A1(n18983), .A2(img[1933]), .B1(n17383), .B2(img[1805]), 
        .O(n16573) );
  AOI22S U19388 ( .A1(n17254), .A2(img[1165]), .B1(n19271), .B2(img[1037]), 
        .O(n16572) );
  AOI22S U19389 ( .A1(n19215), .A2(img[1677]), .B1(n17550), .B2(img[1549]), 
        .O(n16571) );
  AN4S U19390 ( .I1(n16574), .I2(n16573), .I3(n16572), .I4(n16571), .O(n16575)
         );
  AOI22S U19391 ( .A1(n13876), .A2(img[445]), .B1(n13858), .B2(img[317]), .O(
        n16580) );
  AOI22S U19392 ( .A1(n19956), .A2(img[957]), .B1(n13893), .B2(img[829]), .O(
        n16579) );
  AOI22S U19393 ( .A1(n13800), .A2(img[189]), .B1(n17376), .B2(img[61]), .O(
        n16578) );
  AOI22S U19394 ( .A1(n19326), .A2(img[701]), .B1(n13797), .B2(img[573]), .O(
        n16577) );
  AN4S U19395 ( .I1(n16580), .I2(n16579), .I3(n16578), .I4(n16577), .O(n16586)
         );
  AOI22S U19396 ( .A1(n20109), .A2(img[1469]), .B1(n13798), .B2(img[1341]), 
        .O(n16584) );
  AOI22S U19397 ( .A1(n13801), .A2(img[1981]), .B1(n17383), .B2(img[1853]), 
        .O(n16583) );
  AOI22S U19398 ( .A1(n17312), .A2(img[1213]), .B1(n19647), .B2(img[1085]), 
        .O(n16582) );
  AOI22S U19399 ( .A1(n19023), .A2(img[1725]), .B1(n18201), .B2(img[1597]), 
        .O(n16581) );
  AN4S U19400 ( .I1(n16584), .I2(n16583), .I3(n16582), .I4(n16581), .O(n16585)
         );
  AOI22S U19401 ( .A1(n20555), .A2(n13830), .B1(n17928), .B2(n20559), .O(
        n16587) );
  AOI22S U19402 ( .A1(n15506), .A2(img[461]), .B1(n13855), .B2(img[333]), .O(
        n16594) );
  AOI22S U19403 ( .A1(n18946), .A2(img[973]), .B1(n13861), .B2(img[845]), .O(
        n16593) );
  AOI22S U19404 ( .A1(n17354), .A2(img[205]), .B1(n17376), .B2(img[77]), .O(
        n16592) );
  AOI22S U19405 ( .A1(n19641), .A2(img[717]), .B1(n13898), .B2(img[589]), .O(
        n16591) );
  AOI22S U19406 ( .A1(n17382), .A2(img[1485]), .B1(n13798), .B2(img[1357]), 
        .O(n16598) );
  AOI22S U19407 ( .A1(n13841), .A2(img[1997]), .B1(n17383), .B2(img[1869]), 
        .O(n16597) );
  AOI22S U19408 ( .A1(n17347), .A2(img[1229]), .B1(n18922), .B2(img[1101]), 
        .O(n16596) );
  AOI22S U19409 ( .A1(n13867), .A2(img[1741]), .B1(n18201), .B2(img[1613]), 
        .O(n16595) );
  AN4S U19410 ( .I1(n16598), .I2(n16597), .I3(n16596), .I4(n16595), .O(n16599)
         );
  AOI22S U19411 ( .A1(n20032), .A2(img[389]), .B1(n13858), .B2(img[261]), .O(
        n16604) );
  AOI22S U19412 ( .A1(n17810), .A2(img[901]), .B1(n13890), .B2(img[773]), .O(
        n16603) );
  AOI22S U19413 ( .A1(n17330), .A2(img[133]), .B1(n17376), .B2(img[5]), .O(
        n16602) );
  AOI22S U19414 ( .A1(n13875), .A2(img[645]), .B1(n13837), .B2(img[517]), .O(
        n16601) );
  AN4S U19415 ( .I1(n16604), .I2(n16603), .I3(n16602), .I4(n16601), .O(n16610)
         );
  AOI22S U19416 ( .A1(n13823), .A2(img[1413]), .B1(n19182), .B2(img[1285]), 
        .O(n16608) );
  AOI22S U19417 ( .A1(n17793), .A2(img[1925]), .B1(n17617), .B2(img[1797]), 
        .O(n16607) );
  AOI22S U19418 ( .A1(n17254), .A2(img[1157]), .B1(n18922), .B2(img[1029]), 
        .O(n16606) );
  AOI22S U19419 ( .A1(n13786), .A2(img[1669]), .B1(n13796), .B2(img[1541]), 
        .O(n16605) );
  AN4S U19420 ( .I1(n16608), .I2(n16607), .I3(n16606), .I4(n16605), .O(n16609)
         );
  AOI22S U19421 ( .A1(n20546), .A2(n20263), .B1(n13847), .B2(n20558), .O(
        n16665) );
  AOI22S U19422 ( .A1(n15506), .A2(img[453]), .B1(n13858), .B2(img[325]), .O(
        n16614) );
  AOI22S U19423 ( .A1(n18946), .A2(img[965]), .B1(n15653), .B2(img[837]), .O(
        n16613) );
  AOI22S U19424 ( .A1(n17523), .A2(img[197]), .B1(n17376), .B2(img[69]), .O(
        n16612) );
  AOI22S U19425 ( .A1(n19252), .A2(img[709]), .B1(n13797), .B2(img[581]), .O(
        n16611) );
  AN4S U19426 ( .I1(n16614), .I2(n16613), .I3(n16612), .I4(n16611), .O(n16620)
         );
  AOI22S U19427 ( .A1(n17382), .A2(img[1477]), .B1(n13798), .B2(img[1349]), 
        .O(n16618) );
  AOI22S U19428 ( .A1(n17335), .A2(img[1989]), .B1(n17383), .B2(img[1861]), 
        .O(n16617) );
  AOI22S U19429 ( .A1(n17359), .A2(img[1221]), .B1(n19647), .B2(img[1093]), 
        .O(n16616) );
  AOI22S U19430 ( .A1(n13786), .A2(img[1733]), .B1(n18201), .B2(img[1605]), 
        .O(n16615) );
  AN4S U19431 ( .I1(n16618), .I2(n16617), .I3(n16616), .I4(n16615), .O(n16619)
         );
  ND2S U19432 ( .I1(n20539), .I2(n20580), .O(n16664) );
  AOI22S U19433 ( .A1(n20102), .A2(img[413]), .B1(n13858), .B2(img[285]), .O(
        n16624) );
  AOI22S U19434 ( .A1(n13788), .A2(img[925]), .B1(n16048), .B2(img[797]), .O(
        n16623) );
  AOI22S U19435 ( .A1(n18892), .A2(img[157]), .B1(n17376), .B2(img[29]), .O(
        n16622) );
  AOI22S U19436 ( .A1(n19641), .A2(img[669]), .B1(n13898), .B2(img[541]), .O(
        n16621) );
  AN4S U19437 ( .I1(n16624), .I2(n16623), .I3(n16622), .I4(n16621), .O(n16630)
         );
  AOI22S U19438 ( .A1(n20109), .A2(img[1437]), .B1(n17862), .B2(img[1309]), 
        .O(n16628) );
  AOI22S U19439 ( .A1(n19290), .A2(img[1949]), .B1(n17383), .B2(img[1821]), 
        .O(n16627) );
  AOI22S U19440 ( .A1(n17277), .A2(img[1181]), .B1(n13787), .B2(img[1053]), 
        .O(n16626) );
  AOI22S U19441 ( .A1(n20038), .A2(img[1693]), .B1(n13794), .B2(img[1565]), 
        .O(n16625) );
  AN4S U19442 ( .I1(n16628), .I2(n16627), .I3(n16626), .I4(n16625), .O(n16629)
         );
  ND2P U19443 ( .I1(n16630), .I2(n16629), .O(n20545) );
  AOI22S U19444 ( .A1(n18681), .A2(img[501]), .B1(n18262), .B2(img[373]), .O(
        n16634) );
  AOI22S U19445 ( .A1(n18946), .A2(img[1013]), .B1(n15653), .B2(img[885]), .O(
        n16633) );
  AOI22S U19446 ( .A1(n19266), .A2(img[245]), .B1(n17376), .B2(img[117]), .O(
        n16632) );
  AOI22S U19447 ( .A1(n19288), .A2(img[757]), .B1(n13837), .B2(img[629]), .O(
        n16631) );
  AN4S U19448 ( .I1(n16634), .I2(n16633), .I3(n16632), .I4(n16631), .O(n16641)
         );
  AOI22S U19449 ( .A1(n17382), .A2(img[1525]), .B1(n17862), .B2(img[1397]), 
        .O(n16639) );
  AOI22S U19450 ( .A1(n19411), .A2(img[2037]), .B1(n17383), .B2(img[1909]), 
        .O(n16638) );
  AOI22S U19451 ( .A1(n16635), .A2(img[1269]), .B1(n20198), .B2(img[1141]), 
        .O(n16637) );
  AOI22S U19452 ( .A1(n20038), .A2(img[1781]), .B1(n17550), .B2(img[1653]), 
        .O(n16636) );
  AN4S U19453 ( .I1(n16639), .I2(n16638), .I3(n16637), .I4(n16636), .O(n16640)
         );
  AOI22S U19454 ( .A1(n20545), .A2(n13804), .B1(n13846), .B2(n20013), .O(
        n16663) );
  AOI22S U19455 ( .A1(n13876), .A2(img[477]), .B1(n13855), .B2(img[349]), .O(
        n16645) );
  AOI22S U19456 ( .A1(n14505), .A2(img[989]), .B1(n13893), .B2(img[861]), .O(
        n16644) );
  AOI22S U19457 ( .A1(n17218), .A2(img[221]), .B1(n17376), .B2(img[93]), .O(
        n16643) );
  AOI22S U19458 ( .A1(n15568), .A2(img[733]), .B1(n13797), .B2(img[605]), .O(
        n16642) );
  AOI22S U19459 ( .A1(n17382), .A2(img[1501]), .B1(n13798), .B2(img[1373]), 
        .O(n16649) );
  AOI22S U19460 ( .A1(n19411), .A2(img[2013]), .B1(n17383), .B2(img[1885]), 
        .O(n16648) );
  AOI22S U19461 ( .A1(n17347), .A2(img[1245]), .B1(n18548), .B2(img[1117]), 
        .O(n16647) );
  AOI22S U19462 ( .A1(n13863), .A2(img[1757]), .B1(n18201), .B2(img[1629]), 
        .O(n16646) );
  AN4S U19463 ( .I1(n16649), .I2(n16648), .I3(n16647), .I4(n16646), .O(n16650)
         );
  AOI22S U19464 ( .A1(n20102), .A2(img[469]), .B1(n13855), .B2(img[341]), .O(
        n16655) );
  AOI22S U19465 ( .A1(n14822), .A2(img[981]), .B1(n13890), .B2(img[853]), .O(
        n16654) );
  AOI22S U19466 ( .A1(n17218), .A2(img[213]), .B1(n17376), .B2(img[85]), .O(
        n16653) );
  AOI22S U19467 ( .A1(n15568), .A2(img[725]), .B1(n13837), .B2(img[597]), .O(
        n16652) );
  AN4S U19468 ( .I1(n16655), .I2(n16654), .I3(n16653), .I4(n16652), .O(n16661)
         );
  AOI22S U19469 ( .A1(n17382), .A2(img[1493]), .B1(n13798), .B2(img[1365]), 
        .O(n16659) );
  AOI22S U19470 ( .A1(n18773), .A2(img[2005]), .B1(n17383), .B2(img[1877]), 
        .O(n16658) );
  AOI22S U19471 ( .A1(n17277), .A2(img[1237]), .B1(n18548), .B2(img[1109]), 
        .O(n16657) );
  AOI22S U19472 ( .A1(n19215), .A2(img[1749]), .B1(n19715), .B2(img[1621]), 
        .O(n16656) );
  AN4S U19473 ( .I1(n16659), .I2(n16658), .I3(n16657), .I4(n16656), .O(n16660)
         );
  ND2P U19474 ( .I1(n16661), .I2(n16660), .O(n20540) );
  AOI22S U19475 ( .A1(n20561), .A2(n13835), .B1(n13791), .B2(n20540), .O(
        n16662) );
  AN4S U19476 ( .I1(n16665), .I2(n16664), .I3(n16663), .I4(n16662), .O(n16666)
         );
  ND2S U19477 ( .I1(n16667), .I2(n16666), .O(n16704) );
  AOI22S U19478 ( .A1(n16704), .A2(n20364), .B1(n20314), .B2(n16704), .O(
        n16693) );
  AOI22S U19479 ( .A1(n15657), .A2(img[509]), .B1(n13858), .B2(img[381]), .O(
        n16671) );
  AOI22S U19480 ( .A1(n17880), .A2(img[253]), .B1(n19642), .B2(img[125]), .O(
        n16670) );
  AOI22S U19481 ( .A1(n19956), .A2(img[1021]), .B1(n13889), .B2(img[893]), .O(
        n16669) );
  AOI22S U19482 ( .A1(n13886), .A2(img[765]), .B1(n13898), .B2(img[637]), .O(
        n16668) );
  AN4S U19483 ( .I1(n16671), .I2(n16670), .I3(n16669), .I4(n16668), .O(n16677)
         );
  AOI22S U19484 ( .A1(n18910), .A2(img[1277]), .B1(n17885), .B2(img[1149]), 
        .O(n16675) );
  AOI22S U19485 ( .A1(n16075), .A2(img[1789]), .B1(n13796), .B2(img[1661]), 
        .O(n16674) );
  AOI22S U19486 ( .A1(n13823), .A2(img[1533]), .B1(n19001), .B2(img[1405]), 
        .O(n16673) );
  AOI22S U19487 ( .A1(n19411), .A2(img[2045]), .B1(n22928), .B2(img[1917]), 
        .O(n16672) );
  AN4S U19488 ( .I1(n16675), .I2(n16674), .I3(n16673), .I4(n16672), .O(n16676)
         );
  AOI22S U19489 ( .A1(n19603), .A2(n21245), .B1(n20541), .B2(n22923), .O(
        n16679) );
  ND2S U19490 ( .I1(n20541), .I2(n19818), .O(n16678) );
  ND2S U19491 ( .I1(n16679), .I2(n16678), .O(n16680) );
  AOI12HS U19492 ( .B1(n16704), .B2(n19533), .A1(n16680), .O(n16692) );
  BUF1 U19493 ( .I(n18040), .O(n20560) );
  AOI22S U19494 ( .A1(n20558), .A2(n13847), .B1(n20560), .B2(n20539), .O(
        n16684) );
  ND2S U19495 ( .I1(n20557), .I2(n20124), .O(n16683) );
  AOI22S U19496 ( .A1(n20544), .A2(n13839), .B1(n21062), .B2(n20542), .O(
        n16682) );
  AOI22S U19497 ( .A1(n20555), .A2(n13830), .B1(n17938), .B2(n20540), .O(
        n16681) );
  AN4S U19498 ( .I1(n16684), .I2(n16683), .I3(n16682), .I4(n16681), .O(n16690)
         );
  AOI22S U19499 ( .A1(n20551), .A2(n20963), .B1(n17928), .B2(n20559), .O(
        n16688) );
  AOI22S U19500 ( .A1(n20545), .A2(n13804), .B1(n20439), .B2(n20546), .O(
        n16687) );
  AOI22S U19501 ( .A1(n20552), .A2(n17762), .B1(n13846), .B2(n20013), .O(
        n16686) );
  AOI22S U19502 ( .A1(n20543), .A2(n17875), .B1(n13835), .B2(n20561), .O(
        n16685) );
  AN4S U19503 ( .I1(n16688), .I2(n16687), .I3(n16686), .I4(n16685), .O(n16689)
         );
  ND2S U19504 ( .I1(n16690), .I2(n16689), .O(n16740) );
  ND3P U19505 ( .I1(n16693), .I2(n16692), .I3(n16691), .O(n21805) );
  AOI22S U19506 ( .A1(n20542), .A2(n13839), .B1(n17875), .B2(n20557), .O(
        n16697) );
  AOI22S U19507 ( .A1(n20561), .A2(n19483), .B1(n20187), .B2(n20543), .O(
        n16696) );
  AOI22S U19508 ( .A1(n20545), .A2(n20613), .B1(n17762), .B2(n20555), .O(
        n16695) );
  AOI22S U19509 ( .A1(n20558), .A2(n13830), .B1(n17928), .B2(n20551), .O(
        n16694) );
  AN4S U19510 ( .I1(n16697), .I2(n16696), .I3(n16695), .I4(n16694), .O(n16703)
         );
  AOI22S U19511 ( .A1(n20539), .A2(n20439), .B1(n13847), .B2(n20541), .O(
        n16701) );
  ND2S U19512 ( .I1(n20559), .I2(n20524), .O(n16700) );
  AOI22S U19513 ( .A1(n20544), .A2(n13846), .B1(n20438), .B2(n20552), .O(
        n16699) );
  AOI22S U19514 ( .A1(n20546), .A2(n13791), .B1(n19914), .B2(n20540), .O(
        n16698) );
  AN4S U19515 ( .I1(n16701), .I2(n16700), .I3(n16699), .I4(n16698), .O(n16702)
         );
  ND2S U19516 ( .I1(n16703), .I2(n16702), .O(n16739) );
  AOI22S U19517 ( .A1(n16739), .A2(n20364), .B1(n20223), .B2(n16704), .O(
        n16743) );
  AOI22S U19518 ( .A1(n19818), .A2(n20013), .B1(n20013), .B2(n22923), .O(
        n16737) );
  MOAI1 U19519 ( .A1(n16706), .A2(n15142), .B1(n16705), .B2(n13847), .O(n16710) );
  MOAI1 U19520 ( .A1(n16708), .A2(n15448), .B1(n16707), .B2(n13846), .O(n16709) );
  NR2 U19521 ( .I1(n16710), .I2(n16709), .O(n16718) );
  AOI22S U19522 ( .A1(n16712), .A2(n13830), .B1(n20629), .B2(n16711), .O(
        n16717) );
  INV1S U19523 ( .I(n16713), .O(n16714) );
  AOI22S U19524 ( .A1(n16715), .A2(n17762), .B1(n17928), .B2(n16714), .O(
        n16716) );
  ND3 U19525 ( .I1(n16718), .I2(n16717), .I3(n16716), .O(n16735) );
  MOAI1 U19526 ( .A1(n16722), .A2(n13844), .B1(n16721), .B2(n20406), .O(n16723) );
  NR2 U19527 ( .I1(n16724), .I2(n16723), .O(n16733) );
  INV1S U19528 ( .I(n16725), .O(n16726) );
  AOI22S U19529 ( .A1(n16727), .A2(n20439), .B1(n20613), .B2(n16726), .O(
        n16732) );
  INV1S U19530 ( .I(n16728), .O(n16730) );
  AOI22S U19531 ( .A1(n16730), .A2(n17875), .B1(n13839), .B2(n16729), .O(
        n16731) );
  ND3 U19532 ( .I1(n16733), .I2(n16732), .I3(n16731), .O(n16734) );
  NR2P U19533 ( .I1(n16735), .I2(n16734), .O(n20396) );
  INV2 U19534 ( .I(n20396), .O(n20688) );
  AOI22S U19535 ( .A1(n20252), .A2(n21245), .B1(n17686), .B2(n20688), .O(
        n16736) );
  ND2S U19536 ( .I1(n16737), .I2(n16736), .O(n16738) );
  AOI12HS U19537 ( .B1(n16739), .B2(n19533), .A1(n16738), .O(n16742) );
  AN2 U19538 ( .I1(n19608), .I2(n20809), .O(n20062) );
  ND2S U19539 ( .I1(n16740), .I2(n20062), .O(n16741) );
  ND3HT U19540 ( .I1(n16743), .I2(n16742), .I3(n16741), .O(n22055) );
  OAI22S U19541 ( .A1(n29503), .A2(n22054), .B1(n21595), .B2(n22055), .O(
        n17967) );
  ND2P U19542 ( .I1(n22055), .I2(n20809), .O(n21412) );
  INV1S U19543 ( .I(n21412), .O(n21601) );
  AOI22S U19544 ( .A1(n13785), .A2(img[489]), .B1(n19709), .B2(img[361]), .O(
        n16747) );
  AOI22S U19545 ( .A1(n14822), .A2(img[1001]), .B1(n13893), .B2(img[873]), .O(
        n16746) );
  AOI22S U19546 ( .A1(n17729), .A2(img[233]), .B1(n17611), .B2(img[105]), .O(
        n16745) );
  AOI22S U19547 ( .A1(n17730), .A2(img[745]), .B1(n13837), .B2(img[617]), .O(
        n16744) );
  AOI22S U19548 ( .A1(n19193), .A2(img[1513]), .B1(n17862), .B2(img[1385]), 
        .O(n16751) );
  AOI22S U19549 ( .A1(n17778), .A2(img[2025]), .B1(n17863), .B2(img[1897]), 
        .O(n16750) );
  AOI22S U19550 ( .A1(n13827), .A2(img[1257]), .B1(n13802), .B2(img[1129]), 
        .O(n16749) );
  AOI22S U19551 ( .A1(n13786), .A2(img[1769]), .B1(n13794), .B2(img[1641]), 
        .O(n16748) );
  AOI22S U19552 ( .A1(n13883), .A2(img[425]), .B1(n13879), .B2(img[297]), .O(
        n16757) );
  AOI22S U19553 ( .A1(n14822), .A2(img[937]), .B1(n13893), .B2(img[809]), .O(
        n16756) );
  AOI22S U19554 ( .A1(n17249), .A2(img[169]), .B1(n13836), .B2(img[41]), .O(
        n16755) );
  AOI22S U19555 ( .A1(n19326), .A2(img[681]), .B1(n13797), .B2(img[553]), .O(
        n16754) );
  AOI22S U19556 ( .A1(n13823), .A2(img[1449]), .B1(n17862), .B2(img[1321]), 
        .O(n16762) );
  AOI22S U19557 ( .A1(n18819), .A2(img[1961]), .B1(n17863), .B2(img[1833]), 
        .O(n16761) );
  AOI22S U19558 ( .A1(n13783), .A2(img[1193]), .B1(n17712), .B2(img[1065]), 
        .O(n16760) );
  AOI22S U19559 ( .A1(n13867), .A2(img[1705]), .B1(n13796), .B2(img[1577]), 
        .O(n16759) );
  AOI22S U19560 ( .A1(n20444), .A2(n13839), .B1(n17875), .B2(n20445), .O(
        n16829) );
  AOI22S U19561 ( .A1(n20102), .A2(img[433]), .B1(n13896), .B2(img[305]), .O(
        n16768) );
  AOI22S U19562 ( .A1(n19956), .A2(img[945]), .B1(n13889), .B2(img[817]), .O(
        n16767) );
  AOI22S U19563 ( .A1(n19266), .A2(img[177]), .B1(n13836), .B2(img[49]), .O(
        n16766) );
  AOI22S U19564 ( .A1(n13875), .A2(img[689]), .B1(n13898), .B2(img[561]), .O(
        n16765) );
  AOI22S U19565 ( .A1(n19193), .A2(img[1457]), .B1(n13798), .B2(img[1329]), 
        .O(n16772) );
  AOI22S U19566 ( .A1(n18983), .A2(img[1969]), .B1(n17863), .B2(img[1841]), 
        .O(n16771) );
  AOI22S U19567 ( .A1(n13783), .A2(img[1201]), .B1(n17712), .B2(img[1073]), 
        .O(n16770) );
  AOI22S U19568 ( .A1(n19036), .A2(img[1713]), .B1(n13796), .B2(img[1585]), 
        .O(n16769) );
  AOI22S U19569 ( .A1(n13883), .A2(img[481]), .B1(n13896), .B2(img[353]), .O(
        n16778) );
  AOI22S U19570 ( .A1(n18946), .A2(img[993]), .B1(n13893), .B2(img[865]), .O(
        n16777) );
  AOI22S U19571 ( .A1(n17729), .A2(img[225]), .B1(n17611), .B2(img[97]), .O(
        n16776) );
  AOI22S U19572 ( .A1(n17730), .A2(img[737]), .B1(n13837), .B2(img[609]), .O(
        n16775) );
  AOI22S U19573 ( .A1(n19193), .A2(img[1505]), .B1(n17862), .B2(img[1377]), 
        .O(n16782) );
  AOI22S U19574 ( .A1(n20104), .A2(img[2017]), .B1(n17863), .B2(img[1889]), 
        .O(n16781) );
  AOI22S U19575 ( .A1(n14392), .A2(img[1249]), .B1(n13802), .B2(img[1121]), 
        .O(n16780) );
  AOI22S U19576 ( .A1(n19036), .A2(img[1761]), .B1(n13794), .B2(img[1633]), 
        .O(n16779) );
  AOI22S U19577 ( .A1(n20457), .A2(n20187), .B1(n21062), .B2(n20443), .O(
        n16828) );
  AOI22S U19578 ( .A1(n19343), .A2(img[417]), .B1(n13859), .B2(img[289]), .O(
        n16788) );
  AOI22S U19579 ( .A1(n13788), .A2(img[929]), .B1(n13893), .B2(img[801]), .O(
        n16787) );
  AOI22S U19580 ( .A1(n18892), .A2(img[161]), .B1(n20103), .B2(img[33]), .O(
        n16786) );
  AOI22S U19581 ( .A1(n19641), .A2(img[673]), .B1(n13837), .B2(img[545]), .O(
        n16785) );
  AN4S U19582 ( .I1(n16788), .I2(n16787), .I3(n16786), .I4(n16785), .O(n16794)
         );
  AOI22S U19583 ( .A1(n19193), .A2(img[1441]), .B1(n13798), .B2(img[1313]), 
        .O(n16792) );
  AOI22S U19584 ( .A1(n13803), .A2(img[1953]), .B1(n17863), .B2(img[1825]), 
        .O(n16791) );
  AOI22S U19585 ( .A1(n16799), .A2(img[1185]), .B1(n17745), .B2(img[1057]), 
        .O(n16790) );
  AOI22S U19586 ( .A1(n13863), .A2(img[1697]), .B1(n13796), .B2(img[1569]), 
        .O(n16789) );
  AOI22S U19587 ( .A1(n20032), .A2(img[401]), .B1(n13896), .B2(img[273]), .O(
        n16798) );
  AOI22S U19588 ( .A1(n18988), .A2(img[913]), .B1(n13861), .B2(img[785]), .O(
        n16797) );
  AOI22S U19589 ( .A1(n13800), .A2(img[145]), .B1(n17376), .B2(img[17]), .O(
        n16796) );
  AOI22S U19590 ( .A1(n19641), .A2(img[657]), .B1(n13837), .B2(img[529]), .O(
        n16795) );
  AN4S U19591 ( .I1(n16798), .I2(n16797), .I3(n16796), .I4(n16795), .O(n16805)
         );
  AOI22S U19592 ( .A1(n19193), .A2(img[1425]), .B1(n13798), .B2(img[1297]), 
        .O(n16803) );
  AOI22S U19593 ( .A1(n17515), .A2(img[1937]), .B1(n17863), .B2(img[1809]), 
        .O(n16802) );
  AOI22S U19594 ( .A1(n13783), .A2(img[1169]), .B1(n17767), .B2(img[1041]), 
        .O(n16801) );
  AOI22S U19595 ( .A1(n19036), .A2(img[1681]), .B1(n17561), .B2(img[1553]), 
        .O(n16800) );
  AOI22S U19596 ( .A1(n20451), .A2(n20613), .B1(n17762), .B2(n20437), .O(
        n16827) );
  AOI22S U19597 ( .A1(n13825), .A2(img[393]), .B1(n13896), .B2(img[265]), .O(
        n16809) );
  AOI22S U19598 ( .A1(n18946), .A2(img[905]), .B1(n13861), .B2(img[777]), .O(
        n16808) );
  AOI22S U19599 ( .A1(n13800), .A2(img[137]), .B1(n19388), .B2(img[9]), .O(
        n16807) );
  AOI22S U19600 ( .A1(n19252), .A2(img[649]), .B1(n13797), .B2(img[521]), .O(
        n16806) );
  AOI22S U19601 ( .A1(n13803), .A2(img[1929]), .B1(n17863), .B2(img[1801]), 
        .O(n16812) );
  AOI22S U19602 ( .A1(n13827), .A2(img[1161]), .B1(n17767), .B2(img[1033]), 
        .O(n16811) );
  AOI22S U19603 ( .A1(n19023), .A2(img[1673]), .B1(n13794), .B2(img[1545]), 
        .O(n16810) );
  AOI22S U19604 ( .A1(n13883), .A2(img[441]), .B1(n18262), .B2(img[313]), .O(
        n16819) );
  AOI22S U19605 ( .A1(n19649), .A2(img[953]), .B1(n13880), .B2(img[825]), .O(
        n16818) );
  AOI22S U19606 ( .A1(n18713), .A2(img[185]), .B1(n17376), .B2(img[57]), .O(
        n16817) );
  AOI22S U19607 ( .A1(n13875), .A2(img[697]), .B1(n13837), .B2(img[569]), .O(
        n16816) );
  AN4S U19608 ( .I1(n16819), .I2(n16818), .I3(n16817), .I4(n16816), .O(n16825)
         );
  AOI22S U19609 ( .A1(n13823), .A2(img[1465]), .B1(n13798), .B2(img[1337]), 
        .O(n16823) );
  AOI22S U19610 ( .A1(n18983), .A2(img[1977]), .B1(n17863), .B2(img[1849]), 
        .O(n16822) );
  AOI22S U19611 ( .A1(n17277), .A2(img[1209]), .B1(n13802), .B2(img[1081]), 
        .O(n16821) );
  AOI22S U19612 ( .A1(n13867), .A2(img[1721]), .B1(n13794), .B2(img[1593]), 
        .O(n16820) );
  AOI22S U19613 ( .A1(n20456), .A2(n13830), .B1(n17928), .B2(n20455), .O(
        n16826) );
  AN4S U19614 ( .I1(n16829), .I2(n16828), .I3(n16827), .I4(n16826), .O(n16905)
         );
  AOI22S U19615 ( .A1(n13785), .A2(img[457]), .B1(n13879), .B2(img[329]), .O(
        n16833) );
  AOI22S U19616 ( .A1(n16515), .A2(img[969]), .B1(n16048), .B2(img[841]), .O(
        n16832) );
  AOI22S U19617 ( .A1(n17788), .A2(img[201]), .B1(n13836), .B2(img[73]), .O(
        n16831) );
  AOI22S U19618 ( .A1(n16348), .A2(img[713]), .B1(n13797), .B2(img[585]), .O(
        n16830) );
  AOI22S U19619 ( .A1(n13874), .A2(img[1481]), .B1(n17862), .B2(img[1353]), 
        .O(n16837) );
  AOI22S U19620 ( .A1(n18819), .A2(img[1993]), .B1(n17863), .B2(img[1865]), 
        .O(n16836) );
  AOI22S U19621 ( .A1(n17359), .A2(img[1225]), .B1(n13802), .B2(img[1097]), 
        .O(n16835) );
  AOI22S U19622 ( .A1(n16075), .A2(img[1737]), .B1(n13794), .B2(img[1609]), 
        .O(n16834) );
  ND2P U19623 ( .I1(n16839), .I2(n16838), .O(n20446) );
  AOI22S U19624 ( .A1(n20032), .A2(img[385]), .B1(n13858), .B2(img[257]), .O(
        n16843) );
  AOI22S U19625 ( .A1(n18148), .A2(img[897]), .B1(n13861), .B2(img[769]), .O(
        n16842) );
  AOI22S U19626 ( .A1(n17488), .A2(img[129]), .B1(n17611), .B2(img[1]), .O(
        n16841) );
  AOI22S U19627 ( .A1(n19641), .A2(img[641]), .B1(n13797), .B2(img[513]), .O(
        n16840) );
  AN4S U19628 ( .I1(n16843), .I2(n16842), .I3(n16841), .I4(n16840), .O(n16849)
         );
  AOI22S U19629 ( .A1(n13874), .A2(img[1409]), .B1(n13798), .B2(img[1281]), 
        .O(n16847) );
  AOI22S U19630 ( .A1(n17864), .A2(img[1921]), .B1(n17863), .B2(img[1793]), 
        .O(n16846) );
  AOI22S U19631 ( .A1(n17088), .A2(img[1153]), .B1(n13787), .B2(img[1025]), 
        .O(n16845) );
  AOI22S U19632 ( .A1(n19036), .A2(img[1665]), .B1(n17550), .B2(img[1537]), 
        .O(n16844) );
  AOI22S U19633 ( .A1(n20446), .A2(n20263), .B1(n13847), .B2(n20453), .O(
        n16903) );
  AOI22S U19634 ( .A1(n15506), .A2(img[449]), .B1(n13896), .B2(img[321]), .O(
        n16853) );
  AOI22S U19635 ( .A1(n18946), .A2(img[961]), .B1(n13893), .B2(img[833]), .O(
        n16852) );
  AOI22S U19636 ( .A1(n17811), .A2(img[193]), .B1(n17611), .B2(img[65]), .O(
        n16851) );
  AOI22S U19637 ( .A1(n13826), .A2(img[705]), .B1(n13797), .B2(img[577]), .O(
        n16850) );
  AN4S U19638 ( .I1(n16853), .I2(n16852), .I3(n16851), .I4(n16850), .O(n16859)
         );
  AOI22S U19639 ( .A1(n19193), .A2(img[1473]), .B1(n13798), .B2(img[1345]), 
        .O(n16857) );
  AOI22S U19640 ( .A1(n13803), .A2(img[1985]), .B1(n17863), .B2(img[1857]), 
        .O(n16856) );
  AOI22S U19641 ( .A1(n13783), .A2(img[1217]), .B1(n19295), .B2(img[1089]), 
        .O(n16855) );
  AOI22S U19642 ( .A1(n19036), .A2(img[1729]), .B1(n13794), .B2(img[1601]), 
        .O(n16854) );
  ND2S U19643 ( .I1(n20440), .I2(n20580), .O(n16902) );
  AOI22S U19644 ( .A1(n13785), .A2(img[409]), .B1(n19709), .B2(img[281]), .O(
        n16863) );
  AOI22S U19645 ( .A1(n16515), .A2(img[921]), .B1(n13889), .B2(img[793]), .O(
        n16862) );
  AOI22S U19646 ( .A1(n17467), .A2(img[153]), .B1(n17376), .B2(img[25]), .O(
        n16861) );
  AOI22S U19647 ( .A1(n13784), .A2(img[665]), .B1(n13837), .B2(img[537]), .O(
        n16860) );
  AOI22S U19648 ( .A1(n19193), .A2(img[1433]), .B1(n17827), .B2(img[1305]), 
        .O(n16867) );
  AOI22S U19649 ( .A1(n18797), .A2(img[1945]), .B1(n17863), .B2(img[1817]), 
        .O(n16866) );
  AOI22S U19650 ( .A1(n13853), .A2(img[1177]), .B1(n18922), .B2(img[1049]), 
        .O(n16865) );
  AOI22S U19651 ( .A1(n19215), .A2(img[1689]), .B1(n13794), .B2(img[1561]), 
        .O(n16864) );
  AOI22S U19652 ( .A1(n19343), .A2(img[497]), .B1(n13896), .B2(img[369]), .O(
        n16873) );
  AOI22S U19653 ( .A1(n16515), .A2(img[1009]), .B1(n13893), .B2(img[881]), .O(
        n16872) );
  AOI22S U19654 ( .A1(n17330), .A2(img[241]), .B1(n17611), .B2(img[113]), .O(
        n16871) );
  AOI22S U19655 ( .A1(n17835), .A2(img[753]), .B1(n13898), .B2(img[625]), .O(
        n16870) );
  AOI22S U19656 ( .A1(n15630), .A2(img[1521]), .B1(n17862), .B2(img[1393]), 
        .O(n16877) );
  AOI22S U19657 ( .A1(n17793), .A2(img[2033]), .B1(n17863), .B2(img[1905]), 
        .O(n16876) );
  AOI22S U19658 ( .A1(n15315), .A2(img[1265]), .B1(n17840), .B2(img[1137]), 
        .O(n16875) );
  AOI22S U19659 ( .A1(n13867), .A2(img[1777]), .B1(n13794), .B2(img[1649]), 
        .O(n16874) );
  AOI22S U19660 ( .A1(n20452), .A2(n13804), .B1(n13846), .B2(n20458), .O(
        n16901) );
  AOI22S U19661 ( .A1(n13825), .A2(img[473]), .B1(n19709), .B2(img[345]), .O(
        n16883) );
  AOI22S U19662 ( .A1(n20110), .A2(img[985]), .B1(n16048), .B2(img[857]), .O(
        n16882) );
  AOI22S U19663 ( .A1(n17857), .A2(img[217]), .B1(n13836), .B2(img[89]), .O(
        n16881) );
  AOI22S U19664 ( .A1(n19641), .A2(img[729]), .B1(n13837), .B2(img[601]), .O(
        n16880) );
  AOI22S U19665 ( .A1(n13874), .A2(img[1497]), .B1(n17862), .B2(img[1369]), 
        .O(n16887) );
  AOI22S U19666 ( .A1(n13841), .A2(img[2009]), .B1(n17863), .B2(img[1881]), 
        .O(n16886) );
  AOI22S U19667 ( .A1(n17323), .A2(img[1241]), .B1(n17865), .B2(img[1113]), 
        .O(n16885) );
  AOI22S U19668 ( .A1(n13786), .A2(img[1753]), .B1(n13794), .B2(img[1625]), 
        .O(n16884) );
  AOI22S U19669 ( .A1(n13785), .A2(img[465]), .B1(n19709), .B2(img[337]), .O(
        n16893) );
  AOI22S U19670 ( .A1(n18946), .A2(img[977]), .B1(n13893), .B2(img[849]), .O(
        n16892) );
  AOI22S U19671 ( .A1(n17788), .A2(img[209]), .B1(n13836), .B2(img[81]), .O(
        n16891) );
  AOI22S U19672 ( .A1(n16348), .A2(img[721]), .B1(n13797), .B2(img[593]), .O(
        n16890) );
  AOI22S U19673 ( .A1(n19193), .A2(img[1489]), .B1(n17862), .B2(img[1361]), 
        .O(n16897) );
  AOI22S U19674 ( .A1(n13833), .A2(img[2001]), .B1(n17863), .B2(img[1873]), 
        .O(n16896) );
  AOI22S U19675 ( .A1(n17312), .A2(img[1233]), .B1(n17865), .B2(img[1105]), 
        .O(n16895) );
  AOI22S U19676 ( .A1(n18885), .A2(img[1745]), .B1(n13794), .B2(img[1617]), 
        .O(n16894) );
  AN4 U19677 ( .I1(n16897), .I2(n16896), .I3(n16895), .I4(n16894), .O(n16898)
         );
  AOI22S U19678 ( .A1(n20454), .A2(n13835), .B1(n17938), .B2(n20442), .O(
        n16900) );
  AN4S U19679 ( .I1(n16903), .I2(n16902), .I3(n16901), .I4(n16900), .O(n16904)
         );
  AOI22S U19680 ( .A1(n16966), .A2(n20371), .B1(n20364), .B2(n16966), .O(
        n16921) );
  AOI22S U19681 ( .A1(n13825), .A2(img[505]), .B1(n13858), .B2(img[377]), .O(
        n16909) );
  AOI22S U19682 ( .A1(n17880), .A2(img[249]), .B1(n19642), .B2(img[121]), .O(
        n16908) );
  AOI22S U19683 ( .A1(n18946), .A2(img[1017]), .B1(n15653), .B2(img[889]), .O(
        n16907) );
  AOI22S U19684 ( .A1(n13886), .A2(img[761]), .B1(n13837), .B2(img[633]), .O(
        n16906) );
  AN4S U19685 ( .I1(n16909), .I2(n16908), .I3(n16907), .I4(n16906), .O(n16915)
         );
  AOI22S U19686 ( .A1(n18975), .A2(img[1273]), .B1(n17885), .B2(img[1145]), 
        .O(n16913) );
  AOI22S U19687 ( .A1(n13867), .A2(img[1785]), .B1(n18201), .B2(img[1657]), 
        .O(n16912) );
  AOI22S U19688 ( .A1(n17382), .A2(img[1529]), .B1(n19182), .B2(img[1401]), 
        .O(n16911) );
  AOI22S U19689 ( .A1(n13803), .A2(img[2041]), .B1(n22928), .B2(img[1913]), 
        .O(n16910) );
  AOI22S U19690 ( .A1(n19603), .A2(n13887), .B1(n20441), .B2(n22923), .O(
        n16917) );
  ND2S U19691 ( .I1(n20441), .I2(n19818), .O(n16916) );
  ND2S U19692 ( .I1(n16917), .I2(n16916), .O(n16918) );
  AOI12HS U19693 ( .B1(n16966), .B2(n19533), .A1(n16918), .O(n16920) );
  ND2S U19694 ( .I1(n16966), .I2(n19608), .O(n16919) );
  ND3HT U19695 ( .I1(n16921), .I2(n16920), .I3(n16919), .O(n21810) );
  AOI22S U19696 ( .A1(n20443), .A2(n13839), .B1(n17875), .B2(n20451), .O(
        n16925) );
  AOI22S U19697 ( .A1(n20454), .A2(n19483), .B1(n20187), .B2(n20445), .O(
        n16924) );
  AOI22S U19698 ( .A1(n20452), .A2(n20613), .B1(n17762), .B2(n20456), .O(
        n16923) );
  AOI22S U19699 ( .A1(n20453), .A2(n13830), .B1(n17928), .B2(n20457), .O(
        n16922) );
  AN4S U19700 ( .I1(n16925), .I2(n16924), .I3(n16923), .I4(n16922), .O(n16931)
         );
  AOI22S U19701 ( .A1(n20440), .A2(n20439), .B1(n13847), .B2(n20441), .O(
        n16929) );
  ND2S U19702 ( .I1(n20455), .I2(n20524), .O(n16928) );
  AOI22S U19703 ( .A1(n20444), .A2(n13846), .B1(n20438), .B2(n20437), .O(
        n16927) );
  AOI22S U19704 ( .A1(n20446), .A2(n13791), .B1(n13835), .B2(n20442), .O(
        n16926) );
  AN4S U19705 ( .I1(n16929), .I2(n16928), .I3(n16927), .I4(n16926), .O(n16930)
         );
  ND2S U19706 ( .I1(n16931), .I2(n16930), .O(n16965) );
  AOI22S U19707 ( .A1(n16966), .A2(n20223), .B1(n20364), .B2(n16965), .O(
        n16969) );
  AOI22S U19708 ( .A1(n19818), .A2(n20458), .B1(n20458), .B2(n22923), .O(
        n16963) );
  NR2 U19709 ( .I1(n16937), .I2(n16936), .O(n16944) );
  AOI22S U19710 ( .A1(n16939), .A2(n17875), .B1(n20969), .B2(n16938), .O(
        n16943) );
  AOI22S U19711 ( .A1(n16941), .A2(n20613), .B1(n21062), .B2(n16940), .O(
        n16942) );
  ND3 U19712 ( .I1(n16944), .I2(n16943), .I3(n16942), .O(n16961) );
  NR2 U19713 ( .I1(n16950), .I2(n16949), .O(n16959) );
  INV1S U19714 ( .I(n16951), .O(n16952) );
  AOI22S U19715 ( .A1(n16953), .A2(n13830), .B1(n20438), .B2(n16952), .O(
        n16958) );
  INV1S U19716 ( .I(n16954), .O(n16955) );
  AOI22S U19717 ( .A1(n16956), .A2(n13846), .B1(n20629), .B2(n16955), .O(
        n16957) );
  ND3 U19718 ( .I1(n16959), .I2(n16958), .I3(n16957), .O(n16960) );
  NR2T U19719 ( .I1(n16961), .I2(n16960), .O(n20674) );
  INV2 U19720 ( .I(n20674), .O(n20343) );
  AOI22S U19721 ( .A1(n20252), .A2(n13887), .B1(n17686), .B2(n20343), .O(
        n16962) );
  ND2S U19722 ( .I1(n16966), .I2(n20062), .O(n16967) );
  ND3HT U19723 ( .I1(n16969), .I2(n16968), .I3(n16967), .O(n22061) );
  ND2F U19724 ( .I1(n22061), .I2(n20809), .O(n21394) );
  AOI22S U19725 ( .A1(n13883), .A2(img[488]), .B1(n19709), .B2(img[360]), .O(
        n16973) );
  AOI22S U19726 ( .A1(n19037), .A2(img[1000]), .B1(n13890), .B2(img[872]), .O(
        n16972) );
  AOI22S U19727 ( .A1(n17729), .A2(img[232]), .B1(n17611), .B2(img[104]), .O(
        n16971) );
  AOI22S U19728 ( .A1(n17730), .A2(img[744]), .B1(n13797), .B2(img[616]), .O(
        n16970) );
  AN4S U19729 ( .I1(n16973), .I2(n16972), .I3(n16971), .I4(n16970), .O(n16979)
         );
  AOI22S U19730 ( .A1(n13823), .A2(img[1512]), .B1(n17862), .B2(img[1384]), 
        .O(n16977) );
  AOI22S U19731 ( .A1(n17778), .A2(img[2024]), .B1(n17863), .B2(img[1896]), 
        .O(n16976) );
  AOI22S U19732 ( .A1(n14392), .A2(img[1256]), .B1(n13802), .B2(img[1128]), 
        .O(n16975) );
  AOI22S U19733 ( .A1(n19036), .A2(img[1768]), .B1(n13796), .B2(img[1640]), 
        .O(n16974) );
  AN4S U19734 ( .I1(n16977), .I2(n16976), .I3(n16975), .I4(n16974), .O(n16978)
         );
  AOI22S U19735 ( .A1(n13876), .A2(img[424]), .B1(n13858), .B2(img[296]), .O(
        n16983) );
  AOI22S U19736 ( .A1(n14822), .A2(img[936]), .B1(n13893), .B2(img[808]), .O(
        n16982) );
  AOI22S U19737 ( .A1(n19949), .A2(img[168]), .B1(n17611), .B2(img[40]), .O(
        n16981) );
  AOI22S U19738 ( .A1(n13875), .A2(img[680]), .B1(n13837), .B2(img[552]), .O(
        n16980) );
  AN4S U19739 ( .I1(n16983), .I2(n16982), .I3(n16981), .I4(n16980), .O(n16989)
         );
  AOI22S U19740 ( .A1(n13823), .A2(img[1448]), .B1(n19182), .B2(img[1320]), 
        .O(n16987) );
  AOI22S U19741 ( .A1(n13841), .A2(img[1960]), .B1(n17863), .B2(img[1832]), 
        .O(n16986) );
  AOI22S U19742 ( .A1(n13783), .A2(img[1192]), .B1(n17712), .B2(img[1064]), 
        .O(n16985) );
  AOI22S U19743 ( .A1(n13867), .A2(img[1704]), .B1(n13794), .B2(img[1576]), 
        .O(n16984) );
  AOI22S U19744 ( .A1(n21044), .A2(n13839), .B1(n17875), .B2(n21043), .O(
        n17053) );
  AOI22S U19745 ( .A1(n13785), .A2(img[432]), .B1(n13859), .B2(img[304]), .O(
        n16993) );
  AOI22S U19746 ( .A1(n16515), .A2(img[944]), .B1(n15653), .B2(img[816]), .O(
        n16992) );
  AOI22S U19747 ( .A1(n17354), .A2(img[176]), .B1(n19388), .B2(img[48]), .O(
        n16991) );
  AOI22S U19748 ( .A1(n13875), .A2(img[688]), .B1(n13898), .B2(img[560]), .O(
        n16990) );
  AOI22S U19749 ( .A1(n19193), .A2(img[1456]), .B1(n13798), .B2(img[1328]), 
        .O(n16997) );
  AOI22S U19750 ( .A1(n18996), .A2(img[1968]), .B1(n17863), .B2(img[1840]), 
        .O(n16996) );
  AOI22S U19751 ( .A1(n13783), .A2(img[1200]), .B1(n17712), .B2(img[1072]), 
        .O(n16995) );
  AOI22S U19752 ( .A1(n16075), .A2(img[1712]), .B1(n13794), .B2(img[1584]), 
        .O(n16994) );
  AOI22S U19753 ( .A1(n20102), .A2(img[480]), .B1(n13855), .B2(img[352]), .O(
        n17003) );
  AOI22S U19754 ( .A1(n16037), .A2(img[992]), .B1(n15653), .B2(img[864]), .O(
        n17002) );
  AOI22S U19755 ( .A1(n17729), .A2(img[224]), .B1(n17611), .B2(img[96]), .O(
        n17001) );
  AOI22S U19756 ( .A1(n17730), .A2(img[736]), .B1(n13797), .B2(img[608]), .O(
        n17000) );
  AN4S U19757 ( .I1(n17003), .I2(n17002), .I3(n17001), .I4(n17000), .O(n17009)
         );
  AOI22S U19758 ( .A1(n15630), .A2(img[1504]), .B1(n17862), .B2(img[1376]), 
        .O(n17007) );
  AOI22S U19759 ( .A1(n14909), .A2(img[2016]), .B1(n17863), .B2(img[1888]), 
        .O(n17006) );
  AOI22S U19760 ( .A1(n14392), .A2(img[1248]), .B1(n13802), .B2(img[1120]), 
        .O(n17005) );
  AOI22S U19761 ( .A1(n19215), .A2(img[1760]), .B1(n17561), .B2(img[1632]), 
        .O(n17004) );
  AOI22S U19762 ( .A1(n21049), .A2(n20187), .B1(n21062), .B2(n21040), .O(
        n17052) );
  AOI22S U19763 ( .A1(n15506), .A2(img[416]), .B1(n13896), .B2(img[288]), .O(
        n17013) );
  AOI22S U19764 ( .A1(n16515), .A2(img[928]), .B1(n13893), .B2(img[800]), .O(
        n17012) );
  AOI22S U19765 ( .A1(n17600), .A2(img[160]), .B1(n17611), .B2(img[32]), .O(
        n17011) );
  AOI22S U19766 ( .A1(n19641), .A2(img[672]), .B1(n13837), .B2(img[544]), .O(
        n17010) );
  AN4S U19767 ( .I1(n17013), .I2(n17012), .I3(n17011), .I4(n17010), .O(n17019)
         );
  AOI22S U19768 ( .A1(n19193), .A2(img[1440]), .B1(n13798), .B2(img[1312]), 
        .O(n17017) );
  AOI22S U19769 ( .A1(n17515), .A2(img[1952]), .B1(n17863), .B2(img[1824]), 
        .O(n17016) );
  AOI22S U19770 ( .A1(n14392), .A2(img[1184]), .B1(n17745), .B2(img[1056]), 
        .O(n17015) );
  AOI22S U19771 ( .A1(n13786), .A2(img[1696]), .B1(n19416), .B2(img[1568]), 
        .O(n17014) );
  AOI22S U19772 ( .A1(n20032), .A2(img[400]), .B1(n15691), .B2(img[272]), .O(
        n17023) );
  AOI22S U19773 ( .A1(n18946), .A2(img[912]), .B1(n13861), .B2(img[784]), .O(
        n17022) );
  AOI22S U19774 ( .A1(n13800), .A2(img[144]), .B1(n17376), .B2(img[16]), .O(
        n17021) );
  AOI22S U19775 ( .A1(n19641), .A2(img[656]), .B1(n13797), .B2(img[528]), .O(
        n17020) );
  AN4S U19776 ( .I1(n17023), .I2(n17022), .I3(n17021), .I4(n17020), .O(n17029)
         );
  AOI22S U19777 ( .A1(n20109), .A2(img[1424]), .B1(n13798), .B2(img[1296]), 
        .O(n17027) );
  AOI22S U19778 ( .A1(n13801), .A2(img[1936]), .B1(n17863), .B2(img[1808]), 
        .O(n17026) );
  AOI22S U19779 ( .A1(n13783), .A2(img[1168]), .B1(n17767), .B2(img[1040]), 
        .O(n17025) );
  AOI22S U19780 ( .A1(n19036), .A2(img[1680]), .B1(n18201), .B2(img[1552]), 
        .O(n17024) );
  AOI22S U19781 ( .A1(n21058), .A2(n20613), .B1(n17762), .B2(n21050), .O(
        n17051) );
  AOI22S U19782 ( .A1(n13785), .A2(img[392]), .B1(n13859), .B2(img[264]), .O(
        n17033) );
  AOI22S U19783 ( .A1(n16515), .A2(img[904]), .B1(n13890), .B2(img[776]), .O(
        n17032) );
  AOI22S U19784 ( .A1(n13800), .A2(img[136]), .B1(n19388), .B2(img[8]), .O(
        n17031) );
  AOI22S U19785 ( .A1(n19376), .A2(img[648]), .B1(n13837), .B2(img[520]), .O(
        n17030) );
  AN4S U19786 ( .I1(n17033), .I2(n17032), .I3(n17031), .I4(n17030), .O(n17039)
         );
  AOI22S U19787 ( .A1(n19193), .A2(img[1416]), .B1(n17827), .B2(img[1288]), 
        .O(n17037) );
  AOI22S U19788 ( .A1(n13803), .A2(img[1928]), .B1(n17863), .B2(img[1800]), 
        .O(n17036) );
  AOI22S U19789 ( .A1(n13853), .A2(img[1160]), .B1(n17767), .B2(img[1032]), 
        .O(n17035) );
  AOI22S U19790 ( .A1(n19023), .A2(img[1672]), .B1(n18201), .B2(img[1544]), 
        .O(n17034) );
  ND2P U19791 ( .I1(n17039), .I2(n17038), .O(n21054) );
  AOI22S U19792 ( .A1(n19343), .A2(img[440]), .B1(n13896), .B2(img[312]), .O(
        n17043) );
  AOI22S U19793 ( .A1(n13788), .A2(img[952]), .B1(n13890), .B2(img[824]), .O(
        n17042) );
  AOI22S U19794 ( .A1(n17589), .A2(img[184]), .B1(n17611), .B2(img[56]), .O(
        n17041) );
  AOI22S U19795 ( .A1(n13875), .A2(img[696]), .B1(n13898), .B2(img[568]), .O(
        n17040) );
  AN4S U19796 ( .I1(n17043), .I2(n17042), .I3(n17041), .I4(n17040), .O(n17049)
         );
  AOI22S U19797 ( .A1(n13823), .A2(img[1464]), .B1(n13845), .B2(img[1336]), 
        .O(n17047) );
  AOI22S U19798 ( .A1(n18797), .A2(img[1976]), .B1(n17863), .B2(img[1848]), 
        .O(n17046) );
  AOI22S U19799 ( .A1(n15315), .A2(img[1208]), .B1(n13802), .B2(img[1080]), 
        .O(n17045) );
  AOI22S U19800 ( .A1(n13867), .A2(img[1720]), .B1(n13796), .B2(img[1592]), 
        .O(n17044) );
  AN4S U19801 ( .I1(n17047), .I2(n17046), .I3(n17045), .I4(n17044), .O(n17048)
         );
  AOI22S U19802 ( .A1(n21054), .A2(n13830), .B1(n17928), .B2(n21060), .O(
        n17050) );
  AOI22S U19803 ( .A1(n13825), .A2(img[456]), .B1(n13879), .B2(img[328]), .O(
        n17057) );
  AOI22S U19804 ( .A1(n18935), .A2(img[968]), .B1(n16048), .B2(img[840]), .O(
        n17056) );
  AOI22S U19805 ( .A1(n17811), .A2(img[200]), .B1(n19388), .B2(img[72]), .O(
        n17055) );
  AOI22S U19806 ( .A1(n17730), .A2(img[712]), .B1(n13898), .B2(img[584]), .O(
        n17054) );
  AOI22S U19807 ( .A1(n13823), .A2(img[1480]), .B1(n13798), .B2(img[1352]), 
        .O(n17061) );
  AOI22S U19808 ( .A1(n20104), .A2(img[1992]), .B1(n17863), .B2(img[1864]), 
        .O(n17060) );
  AOI22S U19809 ( .A1(n17347), .A2(img[1224]), .B1(n18974), .B2(img[1096]), 
        .O(n17059) );
  AOI22S U19810 ( .A1(n13867), .A2(img[1736]), .B1(n17561), .B2(img[1608]), 
        .O(n17058) );
  ND2P U19811 ( .I1(n17063), .I2(n17062), .O(n21045) );
  AOI22S U19812 ( .A1(n20032), .A2(img[384]), .B1(n13879), .B2(img[256]), .O(
        n17067) );
  AOI22S U19813 ( .A1(n14822), .A2(img[896]), .B1(n13861), .B2(img[768]), .O(
        n17066) );
  AOI22S U19814 ( .A1(n17197), .A2(img[128]), .B1(n17611), .B2(img[0]), .O(
        n17065) );
  AOI22S U19815 ( .A1(n19641), .A2(img[640]), .B1(n13837), .B2(img[512]), .O(
        n17064) );
  AN4S U19816 ( .I1(n17067), .I2(n17066), .I3(n17065), .I4(n17064), .O(n17073)
         );
  AOI22S U19817 ( .A1(n15630), .A2(img[1408]), .B1(n13798), .B2(img[1280]), 
        .O(n17071) );
  AOI22S U19818 ( .A1(n20104), .A2(img[1920]), .B1(n17863), .B2(img[1792]), 
        .O(n17070) );
  AOI22S U19819 ( .A1(n18910), .A2(img[1152]), .B1(n19319), .B2(img[1024]), 
        .O(n17069) );
  AOI22S U19820 ( .A1(n19023), .A2(img[1664]), .B1(n13832), .B2(img[1536]), 
        .O(n17068) );
  AOI22S U19821 ( .A1(n21045), .A2(n20439), .B1(n13847), .B2(n21059), .O(
        n17129) );
  AOI22S U19822 ( .A1(n13883), .A2(img[448]), .B1(n19709), .B2(img[320]), .O(
        n17077) );
  AOI22S U19823 ( .A1(n18148), .A2(img[960]), .B1(n13893), .B2(img[832]), .O(
        n17076) );
  AOI22S U19824 ( .A1(n17811), .A2(img[192]), .B1(n17611), .B2(img[64]), .O(
        n17075) );
  AOI22S U19825 ( .A1(n13875), .A2(img[704]), .B1(n13797), .B2(img[576]), .O(
        n17074) );
  AN4S U19826 ( .I1(n17077), .I2(n17076), .I3(n17075), .I4(n17074), .O(n17083)
         );
  AOI22S U19827 ( .A1(n19193), .A2(img[1472]), .B1(n13798), .B2(img[1344]), 
        .O(n17081) );
  AOI22S U19828 ( .A1(n13801), .A2(img[1984]), .B1(n17863), .B2(img[1856]), 
        .O(n17080) );
  AOI22S U19829 ( .A1(n17088), .A2(img[1216]), .B1(n13792), .B2(img[1088]), 
        .O(n17079) );
  AOI22S U19830 ( .A1(n19036), .A2(img[1728]), .B1(n17550), .B2(img[1600]), 
        .O(n17078) );
  ND2S U19831 ( .I1(n21037), .I2(n20580), .O(n17128) );
  AOI22S U19832 ( .A1(n15657), .A2(img[408]), .B1(n13879), .B2(img[280]), .O(
        n17087) );
  AOI22S U19833 ( .A1(n20110), .A2(img[920]), .B1(n13892), .B2(img[792]), .O(
        n17086) );
  AOI22S U19834 ( .A1(n19266), .A2(img[152]), .B1(n20103), .B2(img[24]), .O(
        n17085) );
  AOI22S U19835 ( .A1(n13784), .A2(img[664]), .B1(n13837), .B2(img[536]), .O(
        n17084) );
  AN4S U19836 ( .I1(n17087), .I2(n17086), .I3(n17085), .I4(n17084), .O(n17094)
         );
  AOI22S U19837 ( .A1(n19193), .A2(img[1432]), .B1(n17827), .B2(img[1304]), 
        .O(n17092) );
  AOI22S U19838 ( .A1(n18773), .A2(img[1944]), .B1(n17863), .B2(img[1816]), 
        .O(n17091) );
  AOI22S U19839 ( .A1(n15315), .A2(img[1176]), .B1(n18922), .B2(img[1048]), 
        .O(n17090) );
  AOI22S U19840 ( .A1(n13786), .A2(img[1688]), .B1(n19715), .B2(img[1560]), 
        .O(n17089) );
  AOI22S U19841 ( .A1(n13785), .A2(img[496]), .B1(n13896), .B2(img[368]), .O(
        n17098) );
  AOI22S U19842 ( .A1(n18935), .A2(img[1008]), .B1(n16048), .B2(img[880]), .O(
        n17097) );
  AOI22S U19843 ( .A1(n19289), .A2(img[240]), .B1(n20103), .B2(img[112]), .O(
        n17096) );
  AOI22S U19844 ( .A1(n17835), .A2(img[752]), .B1(n13797), .B2(img[624]), .O(
        n17095) );
  AN4S U19845 ( .I1(n17098), .I2(n17097), .I3(n17096), .I4(n17095), .O(n17104)
         );
  AOI22S U19846 ( .A1(n15630), .A2(img[1520]), .B1(n17862), .B2(img[1392]), 
        .O(n17102) );
  AOI22S U19847 ( .A1(n18996), .A2(img[2032]), .B1(n17863), .B2(img[1904]), 
        .O(n17101) );
  AOI22S U19848 ( .A1(n16799), .A2(img[1264]), .B1(n17840), .B2(img[1136]), 
        .O(n17100) );
  AOI22S U19849 ( .A1(n19036), .A2(img[1776]), .B1(n17550), .B2(img[1648]), 
        .O(n17099) );
  AOI22S U19850 ( .A1(n21046), .A2(n13804), .B1(n13846), .B2(n21053), .O(
        n17127) );
  AOI22S U19851 ( .A1(n13876), .A2(img[472]), .B1(n19709), .B2(img[344]), .O(
        n17108) );
  AOI22S U19852 ( .A1(n19037), .A2(img[984]), .B1(n16048), .B2(img[856]), .O(
        n17107) );
  AOI22S U19853 ( .A1(n17857), .A2(img[216]), .B1(n17611), .B2(img[88]), .O(
        n17106) );
  AOI22S U19854 ( .A1(n19641), .A2(img[728]), .B1(n13797), .B2(img[600]), .O(
        n17105) );
  AN4S U19855 ( .I1(n17108), .I2(n17107), .I3(n17106), .I4(n17105), .O(n17114)
         );
  AOI22S U19856 ( .A1(n13823), .A2(img[1496]), .B1(n17827), .B2(img[1368]), 
        .O(n17112) );
  AOI22S U19857 ( .A1(n18958), .A2(img[2008]), .B1(n17863), .B2(img[1880]), 
        .O(n17111) );
  AOI22S U19858 ( .A1(n17254), .A2(img[1240]), .B1(n17865), .B2(img[1112]), 
        .O(n17110) );
  AOI22S U19859 ( .A1(n19023), .A2(img[1752]), .B1(n13794), .B2(img[1624]), 
        .O(n17109) );
  AOI22S U19860 ( .A1(n13785), .A2(img[464]), .B1(n13855), .B2(img[336]), .O(
        n17119) );
  AOI22S U19861 ( .A1(n20110), .A2(img[976]), .B1(n13893), .B2(img[848]), .O(
        n17118) );
  AOI22S U19862 ( .A1(n17788), .A2(img[208]), .B1(n17611), .B2(img[80]), .O(
        n17117) );
  AOI22S U19863 ( .A1(n16348), .A2(img[720]), .B1(n13797), .B2(img[592]), .O(
        n17116) );
  AN4S U19864 ( .I1(n17119), .I2(n17118), .I3(n17117), .I4(n17116), .O(n17125)
         );
  AOI22S U19865 ( .A1(n13823), .A2(img[1488]), .B1(n17827), .B2(img[1360]), 
        .O(n17123) );
  AOI22S U19866 ( .A1(n17793), .A2(img[2000]), .B1(n17863), .B2(img[1872]), 
        .O(n17122) );
  AOI22S U19867 ( .A1(n17336), .A2(img[1232]), .B1(n19955), .B2(img[1104]), 
        .O(n17121) );
  AOI22S U19868 ( .A1(n13786), .A2(img[1744]), .B1(n13794), .B2(img[1616]), 
        .O(n17120) );
  AOI22S U19869 ( .A1(n21063), .A2(n19914), .B1(n17938), .B2(n21038), .O(
        n17126) );
  AOI22S U19870 ( .A1(n17191), .A2(n20371), .B1(n20364), .B2(n17191), .O(
        n17147) );
  AOI22S U19871 ( .A1(n13825), .A2(img[504]), .B1(n13858), .B2(img[376]), .O(
        n17135) );
  AOI22S U19872 ( .A1(n17880), .A2(img[248]), .B1(n19642), .B2(img[120]), .O(
        n17134) );
  AOI22S U19873 ( .A1(n20110), .A2(img[1016]), .B1(n13890), .B2(img[888]), .O(
        n17133) );
  AOI22S U19874 ( .A1(n13886), .A2(img[760]), .B1(n13797), .B2(img[632]), .O(
        n17132) );
  AN4S U19875 ( .I1(n17135), .I2(n17134), .I3(n17133), .I4(n17132), .O(n17141)
         );
  AOI22S U19876 ( .A1(n17254), .A2(img[1272]), .B1(n17885), .B2(img[1144]), 
        .O(n17139) );
  AOI22S U19877 ( .A1(n19036), .A2(img[1784]), .B1(n18201), .B2(img[1656]), 
        .O(n17138) );
  AOI22S U19878 ( .A1(n17382), .A2(img[1528]), .B1(n18751), .B2(img[1400]), 
        .O(n17137) );
  AOI22S U19879 ( .A1(n17793), .A2(img[2040]), .B1(n22928), .B2(img[1912]), 
        .O(n17136) );
  AN4S U19880 ( .I1(n17139), .I2(n17138), .I3(n17137), .I4(n17136), .O(n17140)
         );
  ND2P U19881 ( .I1(n17141), .I2(n17140), .O(n21039) );
  AOI22S U19882 ( .A1(n19603), .A2(n20345), .B1(n21039), .B2(n22923), .O(
        n17143) );
  ND2S U19883 ( .I1(n21039), .I2(n19818), .O(n17142) );
  ND2S U19884 ( .I1(n17143), .I2(n17142), .O(n17144) );
  AOI12HS U19885 ( .B1(n17191), .B2(n19533), .A1(n17144), .O(n17146) );
  ND2S U19886 ( .I1(n17191), .I2(n19608), .O(n17145) );
  ND3P U19887 ( .I1(n17147), .I2(n17146), .I3(n17145), .O(n21809) );
  AOI12HS U19888 ( .B1(n22121), .B2(n21810), .A1(n21809), .O(n17196) );
  AOI22S U19889 ( .A1(n21040), .A2(n13839), .B1(n17875), .B2(n21058), .O(
        n17151) );
  AOI22S U19890 ( .A1(n21063), .A2(n19483), .B1(n20187), .B2(n21043), .O(
        n17150) );
  AOI22S U19891 ( .A1(n21046), .A2(n20613), .B1(n17762), .B2(n21054), .O(
        n17149) );
  AOI22S U19892 ( .A1(n21059), .A2(n13830), .B1(n17928), .B2(n21049), .O(
        n17148) );
  AN4S U19893 ( .I1(n17151), .I2(n17150), .I3(n17149), .I4(n17148), .O(n17157)
         );
  AOI22S U19894 ( .A1(n21037), .A2(n20439), .B1(n13847), .B2(n21039), .O(
        n17155) );
  ND2S U19895 ( .I1(n21060), .I2(n20580), .O(n17154) );
  AOI22S U19896 ( .A1(n21044), .A2(n13846), .B1(n20438), .B2(n21050), .O(
        n17153) );
  AOI22S U19897 ( .A1(n21045), .A2(n13791), .B1(n13835), .B2(n21038), .O(
        n17152) );
  AN4S U19898 ( .I1(n17155), .I2(n17154), .I3(n17153), .I4(n17152), .O(n17156)
         );
  ND2S U19899 ( .I1(n17157), .I2(n17156), .O(n17190) );
  AOI22S U19900 ( .A1(n17191), .A2(n20223), .B1(n20364), .B2(n17190), .O(
        n17194) );
  ND2P U19901 ( .I1(n19573), .I2(n20809), .O(n21641) );
  INV1 U19902 ( .I(n21641), .O(n21260) );
  OR2 U19903 ( .I1(n19473), .I2(n19700), .O(n19871) );
  INV2 U19904 ( .I(n19871), .O(n20373) );
  ND2 U19905 ( .I1(n21260), .I2(n20373), .O(n17188) );
  NR2 U19906 ( .I1(n17163), .I2(n17162), .O(n17170) );
  AOI22S U19907 ( .A1(n17167), .A2(n13793), .B1(n17166), .B2(n20969), .O(
        n17168) );
  ND3 U19908 ( .I1(n17170), .I2(n17169), .I3(n17168), .O(n17185) );
  NR2 U19909 ( .I1(n17176), .I2(n17175), .O(n17183) );
  AOI22S U19910 ( .A1(n13839), .A2(n17178), .B1(n17177), .B2(n13847), .O(
        n17182) );
  AOI22S U19911 ( .A1(n17875), .A2(n17180), .B1(n17179), .B2(n13804), .O(
        n17181) );
  ND3 U19912 ( .I1(n17183), .I2(n17182), .I3(n17181), .O(n17184) );
  NR2P U19913 ( .I1(n17185), .I2(n17184), .O(n20386) );
  INV2 U19914 ( .I(n20386), .O(n20977) );
  ND2S U19915 ( .I1(n17686), .I2(n20977), .O(n17187) );
  AOI12HS U19916 ( .B1(n19818), .B2(n21053), .A1(n13943), .O(n17186) );
  ND3 U19917 ( .I1(n17188), .I2(n17187), .I3(n17186), .O(n17189) );
  AOI12HS U19918 ( .B1(n17190), .B2(n19533), .A1(n17189), .O(n17193) );
  ND2S U19919 ( .I1(n17191), .I2(n20062), .O(n17192) );
  ND3P U19920 ( .I1(n17194), .I2(n17193), .I3(n17192), .O(n22060) );
  NR2F U19921 ( .I1(n13822), .I2(n17195), .O(n21643) );
  MOAI1 U19922 ( .A1(n21810), .A2(n21394), .B1(n17196), .B2(n21643), .O(n17697) );
  AOI22S U19923 ( .A1(n20032), .A2(img[482]), .B1(n13858), .B2(img[354]), .O(
        n17201) );
  AOI22S U19924 ( .A1(n14189), .A2(img[994]), .B1(n13893), .B2(img[866]), .O(
        n17200) );
  AOI22S U19925 ( .A1(n17197), .A2(img[226]), .B1(n17376), .B2(img[98]), .O(
        n17199) );
  AOI22S U19926 ( .A1(n19376), .A2(img[738]), .B1(n13797), .B2(img[610]), .O(
        n17198) );
  AN4S U19927 ( .I1(n17201), .I2(n17200), .I3(n17199), .I4(n17198), .O(n17207)
         );
  AOI22S U19928 ( .A1(n17382), .A2(img[1506]), .B1(n13798), .B2(img[1378]), 
        .O(n17205) );
  AOI22S U19929 ( .A1(n17515), .A2(img[2018]), .B1(n17383), .B2(img[1890]), 
        .O(n17204) );
  AOI22S U19930 ( .A1(n15315), .A2(img[1250]), .B1(n18623), .B2(img[1122]), 
        .O(n17203) );
  AOI22S U19931 ( .A1(n19036), .A2(img[1762]), .B1(n18201), .B2(img[1634]), 
        .O(n17202) );
  AN4S U19932 ( .I1(n17205), .I2(n17204), .I3(n17203), .I4(n17202), .O(n17206)
         );
  AOI22S U19933 ( .A1(n20102), .A2(img[418]), .B1(n13858), .B2(img[290]), .O(
        n17211) );
  AOI22S U19934 ( .A1(n14822), .A2(img[930]), .B1(n13893), .B2(img[802]), .O(
        n17210) );
  AOI22S U19935 ( .A1(n17249), .A2(img[162]), .B1(n17376), .B2(img[34]), .O(
        n17209) );
  AOI22S U19936 ( .A1(n13826), .A2(img[674]), .B1(n13898), .B2(img[546]), .O(
        n17208) );
  AN4S U19937 ( .I1(n17211), .I2(n17210), .I3(n17209), .I4(n17208), .O(n17217)
         );
  AOI22S U19938 ( .A1(n19193), .A2(img[1442]), .B1(n13799), .B2(img[1314]), 
        .O(n17215) );
  AOI22S U19939 ( .A1(n18996), .A2(img[1954]), .B1(n17383), .B2(img[1826]), 
        .O(n17214) );
  AOI22S U19940 ( .A1(n17277), .A2(img[1186]), .B1(n13787), .B2(img[1058]), 
        .O(n17213) );
  AOI22S U19941 ( .A1(n19215), .A2(img[1698]), .B1(n17550), .B2(img[1570]), 
        .O(n17212) );
  AN4S U19942 ( .I1(n17215), .I2(n17214), .I3(n17213), .I4(n17212), .O(n17216)
         );
  AOI22S U19943 ( .A1(n20471), .A2(n13839), .B1(n17875), .B2(n20489), .O(
        n17287) );
  AOI22S U19944 ( .A1(n15657), .A2(img[474]), .B1(n13896), .B2(img[346]), .O(
        n17222) );
  AOI22S U19945 ( .A1(n18946), .A2(img[986]), .B1(n13880), .B2(img[858]), .O(
        n17221) );
  AOI22S U19946 ( .A1(n17218), .A2(img[218]), .B1(n17376), .B2(img[90]), .O(
        n17220) );
  AOI22S U19947 ( .A1(n19641), .A2(img[730]), .B1(n13837), .B2(img[602]), .O(
        n17219) );
  AN4S U19948 ( .I1(n17222), .I2(n17221), .I3(n17220), .I4(n17219), .O(n17228)
         );
  AOI22S U19949 ( .A1(n17382), .A2(img[1498]), .B1(n13798), .B2(img[1370]), 
        .O(n17226) );
  AOI22S U19950 ( .A1(n19290), .A2(img[2010]), .B1(n17383), .B2(img[1882]), 
        .O(n17225) );
  AOI22S U19951 ( .A1(n17254), .A2(img[1242]), .B1(n18548), .B2(img[1114]), 
        .O(n17224) );
  AOI22S U19952 ( .A1(n19023), .A2(img[1754]), .B1(n18201), .B2(img[1626]), 
        .O(n17223) );
  AN4S U19953 ( .I1(n17226), .I2(n17225), .I3(n17224), .I4(n17223), .O(n17227)
         );
  AOI22S U19954 ( .A1(n13785), .A2(img[426]), .B1(n13858), .B2(img[298]), .O(
        n17232) );
  AOI22S U19955 ( .A1(n18946), .A2(img[938]), .B1(n13861), .B2(img[810]), .O(
        n17231) );
  AOI22S U19956 ( .A1(n17271), .A2(img[170]), .B1(n17376), .B2(img[42]), .O(
        n17230) );
  AOI22S U19957 ( .A1(n17730), .A2(img[682]), .B1(n13797), .B2(img[554]), .O(
        n17229) );
  AN4S U19958 ( .I1(n17232), .I2(n17231), .I3(n17230), .I4(n17229), .O(n17238)
         );
  AOI22S U19959 ( .A1(n20109), .A2(img[1450]), .B1(n17827), .B2(img[1322]), 
        .O(n17236) );
  AOI22S U19960 ( .A1(n14909), .A2(img[1962]), .B1(n17383), .B2(img[1834]), 
        .O(n17235) );
  AOI22S U19961 ( .A1(n17312), .A2(img[1194]), .B1(n17276), .B2(img[1066]), 
        .O(n17234) );
  AOI22S U19962 ( .A1(n19215), .A2(img[1706]), .B1(n18201), .B2(img[1578]), 
        .O(n17233) );
  AN4S U19963 ( .I1(n17236), .I2(n17235), .I3(n17234), .I4(n17233), .O(n17237)
         );
  ND2P U19964 ( .I1(n17238), .I2(n17237), .O(n20474) );
  AOI22S U19965 ( .A1(n20492), .A2(n19483), .B1(n20187), .B2(n20474), .O(
        n17286) );
  AOI22S U19966 ( .A1(n15506), .A2(img[410]), .B1(n19709), .B2(img[282]), .O(
        n17242) );
  AOI22S U19967 ( .A1(n16515), .A2(img[922]), .B1(n13890), .B2(img[794]), .O(
        n17241) );
  AOI22S U19968 ( .A1(n17330), .A2(img[154]), .B1(n17376), .B2(img[26]), .O(
        n17240) );
  AOI22S U19969 ( .A1(n19641), .A2(img[666]), .B1(n13797), .B2(img[538]), .O(
        n17239) );
  AN4S U19970 ( .I1(n17242), .I2(n17241), .I3(n17240), .I4(n17239), .O(n17248)
         );
  AOI22S U19971 ( .A1(n13823), .A2(img[1434]), .B1(n17827), .B2(img[1306]), 
        .O(n17246) );
  AOI22S U19972 ( .A1(n17515), .A2(img[1946]), .B1(n17383), .B2(img[1818]), 
        .O(n17245) );
  AOI22S U19973 ( .A1(n17254), .A2(img[1178]), .B1(n18922), .B2(img[1050]), 
        .O(n17244) );
  AOI22S U19974 ( .A1(n19036), .A2(img[1690]), .B1(n18201), .B2(img[1562]), 
        .O(n17243) );
  AN4S U19975 ( .I1(n17246), .I2(n17245), .I3(n17244), .I4(n17243), .O(n17247)
         );
  AOI22S U19976 ( .A1(n19343), .A2(img[394]), .B1(n13855), .B2(img[266]), .O(
        n17253) );
  AOI22S U19977 ( .A1(n18911), .A2(img[906]), .B1(n16048), .B2(img[778]), .O(
        n17252) );
  AOI22S U19978 ( .A1(n17249), .A2(img[138]), .B1(n17376), .B2(img[10]), .O(
        n17251) );
  AOI22S U19979 ( .A1(n18702), .A2(img[650]), .B1(n13797), .B2(img[522]), .O(
        n17250) );
  AN4S U19980 ( .I1(n17253), .I2(n17252), .I3(n17251), .I4(n17250), .O(n17260)
         );
  AOI22S U19981 ( .A1(n19193), .A2(img[1418]), .B1(n13845), .B2(img[1290]), 
        .O(n17258) );
  AOI22S U19982 ( .A1(n13801), .A2(img[1930]), .B1(n17383), .B2(img[1802]), 
        .O(n17257) );
  AOI22S U19983 ( .A1(n17254), .A2(img[1162]), .B1(n17767), .B2(img[1034]), 
        .O(n17256) );
  AOI22S U19984 ( .A1(n19023), .A2(img[1674]), .B1(n17561), .B2(img[1546]), 
        .O(n17255) );
  AN4S U19985 ( .I1(n17258), .I2(n17257), .I3(n17256), .I4(n17255), .O(n17259)
         );
  AOI22S U19986 ( .A1(n20477), .A2(n20613), .B1(n17762), .B2(n20485), .O(
        n17285) );
  AOI22S U19987 ( .A1(n20032), .A2(img[386]), .B1(n13855), .B2(img[258]), .O(
        n17264) );
  AOI22S U19988 ( .A1(n18935), .A2(img[898]), .B1(n13880), .B2(img[770]), .O(
        n17263) );
  AOI22S U19989 ( .A1(n17218), .A2(img[130]), .B1(n17376), .B2(img[2]), .O(
        n17262) );
  AOI22S U19990 ( .A1(n17835), .A2(img[642]), .B1(n13837), .B2(img[514]), .O(
        n17261) );
  AN4S U19991 ( .I1(n17264), .I2(n17263), .I3(n17262), .I4(n17261), .O(n17270)
         );
  AOI22S U19992 ( .A1(n13823), .A2(img[1410]), .B1(n13845), .B2(img[1282]), 
        .O(n17268) );
  AOI22S U19993 ( .A1(n18797), .A2(img[1922]), .B1(n19950), .B2(img[1794]), 
        .O(n17267) );
  AOI22S U19994 ( .A1(n17323), .A2(img[1154]), .B1(n18922), .B2(img[1026]), 
        .O(n17266) );
  AOI22S U19995 ( .A1(n19215), .A2(img[1666]), .B1(n13794), .B2(img[1538]), 
        .O(n17265) );
  AN4S U19996 ( .I1(n17268), .I2(n17267), .I3(n17266), .I4(n17265), .O(n17269)
         );
  AOI22S U19997 ( .A1(n20102), .A2(img[434]), .B1(n13859), .B2(img[306]), .O(
        n17275) );
  AOI22S U19998 ( .A1(n18946), .A2(img[946]), .B1(n13893), .B2(img[818]), .O(
        n17274) );
  AOI22S U19999 ( .A1(n17271), .A2(img[178]), .B1(n17376), .B2(img[50]), .O(
        n17273) );
  AOI22S U20000 ( .A1(n19342), .A2(img[690]), .B1(n13837), .B2(img[562]), .O(
        n17272) );
  AN4S U20001 ( .I1(n17275), .I2(n17274), .I3(n17273), .I4(n17272), .O(n17283)
         );
  AOI22S U20002 ( .A1(n20109), .A2(img[1458]), .B1(n13798), .B2(img[1330]), 
        .O(n17281) );
  AOI22S U20003 ( .A1(n13841), .A2(img[1970]), .B1(n17383), .B2(img[1842]), 
        .O(n17280) );
  AOI22S U20004 ( .A1(n17277), .A2(img[1202]), .B1(n17276), .B2(img[1074]), 
        .O(n17279) );
  AOI22S U20005 ( .A1(n19036), .A2(img[1714]), .B1(n19416), .B2(img[1586]), 
        .O(n17278) );
  AN4S U20006 ( .I1(n17281), .I2(n17280), .I3(n17279), .I4(n17278), .O(n17282)
         );
  AOI22S U20007 ( .A1(n20490), .A2(n13830), .B1(n17928), .B2(n20480), .O(
        n17284) );
  AN4S U20008 ( .I1(n17287), .I2(n17286), .I3(n17285), .I4(n17284), .O(n17371)
         );
  AOI22S U20009 ( .A1(n13876), .A2(img[450]), .B1(n13858), .B2(img[322]), .O(
        n17291) );
  AOI22S U20010 ( .A1(n20110), .A2(img[962]), .B1(n13861), .B2(img[834]), .O(
        n17290) );
  AOI22S U20011 ( .A1(n17271), .A2(img[194]), .B1(n17376), .B2(img[66]), .O(
        n17289) );
  AOI22S U20012 ( .A1(n13875), .A2(img[706]), .B1(n13898), .B2(img[578]), .O(
        n17288) );
  AN4S U20013 ( .I1(n17291), .I2(n17290), .I3(n17289), .I4(n17288), .O(n17297)
         );
  AOI22S U20014 ( .A1(n20109), .A2(img[1474]), .B1(n13798), .B2(img[1346]), 
        .O(n17295) );
  AOI22S U20015 ( .A1(n13841), .A2(img[1986]), .B1(n17383), .B2(img[1858]), 
        .O(n17294) );
  AOI22S U20016 ( .A1(n17359), .A2(img[1218]), .B1(n19647), .B2(img[1090]), 
        .O(n17293) );
  AOI22S U20017 ( .A1(n19023), .A2(img[1730]), .B1(n18201), .B2(img[1602]), 
        .O(n17292) );
  AN4S U20018 ( .I1(n17295), .I2(n17294), .I3(n17293), .I4(n17292), .O(n17296)
         );
  AOI22S U20019 ( .A1(n13825), .A2(img[506]), .B1(n13858), .B2(img[378]), .O(
        n17301) );
  AOI22S U20020 ( .A1(n17880), .A2(img[250]), .B1(n19642), .B2(img[122]), .O(
        n17300) );
  AOI22S U20021 ( .A1(n14505), .A2(img[1018]), .B1(n13877), .B2(img[890]), .O(
        n17299) );
  AOI22S U20022 ( .A1(n13886), .A2(img[762]), .B1(n13797), .B2(img[634]), .O(
        n17298) );
  AN4S U20023 ( .I1(n17301), .I2(n17300), .I3(n17299), .I4(n17298), .O(n17307)
         );
  AOI22S U20024 ( .A1(n18897), .A2(img[1274]), .B1(n17885), .B2(img[1146]), 
        .O(n17305) );
  AOI22S U20025 ( .A1(n18885), .A2(img[1786]), .B1(n18201), .B2(img[1658]), 
        .O(n17304) );
  AOI22S U20026 ( .A1(n20109), .A2(img[1530]), .B1(n17862), .B2(img[1402]), 
        .O(n17303) );
  AOI22S U20027 ( .A1(n13841), .A2(img[2042]), .B1(n22928), .B2(img[1914]), 
        .O(n17302) );
  AN4S U20028 ( .I1(n17305), .I2(n17304), .I3(n17303), .I4(n17302), .O(n17306)
         );
  ND2P U20029 ( .I1(n17307), .I2(n17306), .O(n20470) );
  AOI22S U20030 ( .A1(n20468), .A2(n20439), .B1(n13847), .B2(n20470), .O(
        n17369) );
  AOI22S U20031 ( .A1(n13785), .A2(img[442]), .B1(n13858), .B2(img[314]), .O(
        n17311) );
  AOI22S U20032 ( .A1(n18988), .A2(img[954]), .B1(n15653), .B2(img[826]), .O(
        n17310) );
  AOI22S U20033 ( .A1(n17377), .A2(img[186]), .B1(n17376), .B2(img[58]), .O(
        n17309) );
  AOI22S U20034 ( .A1(n19288), .A2(img[698]), .B1(n13898), .B2(img[570]), .O(
        n17308) );
  AN4S U20035 ( .I1(n17311), .I2(n17310), .I3(n17309), .I4(n17308), .O(n17318)
         );
  AOI22S U20036 ( .A1(n20109), .A2(img[1466]), .B1(n13845), .B2(img[1338]), 
        .O(n17316) );
  AOI22S U20037 ( .A1(n17816), .A2(img[1978]), .B1(n17383), .B2(img[1850]), 
        .O(n17315) );
  AOI22S U20038 ( .A1(n17312), .A2(img[1210]), .B1(n19647), .B2(img[1082]), 
        .O(n17314) );
  AOI22S U20039 ( .A1(n19215), .A2(img[1722]), .B1(n18201), .B2(img[1594]), 
        .O(n17313) );
  AN4S U20040 ( .I1(n17316), .I2(n17315), .I3(n17314), .I4(n17313), .O(n17317)
         );
  ND2P U20041 ( .I1(n17318), .I2(n17317), .O(n20491) );
  ND2S U20042 ( .I1(n20491), .I2(n20524), .O(n17368) );
  AOI22S U20043 ( .A1(n13825), .A2(img[490]), .B1(n13858), .B2(img[362]), .O(
        n17322) );
  AOI22S U20044 ( .A1(n14505), .A2(img[1002]), .B1(n17115), .B2(img[874]), .O(
        n17321) );
  AOI22S U20045 ( .A1(n17377), .A2(img[234]), .B1(n17376), .B2(img[106]), .O(
        n17320) );
  AOI22S U20046 ( .A1(n19641), .A2(img[746]), .B1(n13898), .B2(img[618]), .O(
        n17319) );
  AN4S U20047 ( .I1(n17322), .I2(n17321), .I3(n17320), .I4(n17319), .O(n17329)
         );
  AOI22S U20048 ( .A1(n17382), .A2(img[1514]), .B1(n19182), .B2(img[1386]), 
        .O(n17327) );
  AOI22S U20049 ( .A1(n13833), .A2(img[2026]), .B1(n17383), .B2(img[1898]), 
        .O(n17326) );
  AOI22S U20050 ( .A1(n17323), .A2(img[1258]), .B1(n13787), .B2(img[1130]), 
        .O(n17325) );
  AOI22S U20051 ( .A1(n15751), .A2(img[1770]), .B1(n18201), .B2(img[1642]), 
        .O(n17324) );
  AN4S U20052 ( .I1(n17327), .I2(n17326), .I3(n17325), .I4(n17324), .O(n17328)
         );
  AOI22S U20053 ( .A1(n13825), .A2(img[402]), .B1(n13858), .B2(img[274]), .O(
        n17334) );
  AOI22S U20054 ( .A1(n16037), .A2(img[914]), .B1(n15653), .B2(img[786]), .O(
        n17333) );
  AOI22S U20055 ( .A1(n17330), .A2(img[146]), .B1(n17376), .B2(img[18]), .O(
        n17332) );
  AOI22S U20056 ( .A1(n19265), .A2(img[658]), .B1(n13797), .B2(img[530]), .O(
        n17331) );
  AN4S U20057 ( .I1(n17334), .I2(n17333), .I3(n17332), .I4(n17331), .O(n17342)
         );
  AOI22S U20058 ( .A1(n19193), .A2(img[1426]), .B1(n17862), .B2(img[1298]), 
        .O(n17340) );
  AOI22S U20059 ( .A1(n13803), .A2(img[1938]), .B1(n17383), .B2(img[1810]), 
        .O(n17339) );
  AOI22S U20060 ( .A1(n17336), .A2(img[1170]), .B1(n18922), .B2(img[1042]), 
        .O(n17338) );
  AOI22S U20061 ( .A1(n19036), .A2(img[1682]), .B1(n13794), .B2(img[1554]), 
        .O(n17337) );
  AN4S U20062 ( .I1(n17340), .I2(n17339), .I3(n17338), .I4(n17337), .O(n17341)
         );
  AOI22S U20063 ( .A1(n20475), .A2(n13846), .B1(n20438), .B2(n20481), .O(
        n17367) );
  AOI22S U20064 ( .A1(n13883), .A2(img[458]), .B1(n13879), .B2(img[330]), .O(
        n17346) );
  AOI22S U20065 ( .A1(n16037), .A2(img[970]), .B1(n15653), .B2(img[842]), .O(
        n17345) );
  AOI22S U20066 ( .A1(n17354), .A2(img[202]), .B1(n17376), .B2(img[74]), .O(
        n17344) );
  AOI22S U20067 ( .A1(n19641), .A2(img[714]), .B1(n13837), .B2(img[586]), .O(
        n17343) );
  AN4S U20068 ( .I1(n17346), .I2(n17345), .I3(n17344), .I4(n17343), .O(n17353)
         );
  AOI22S U20069 ( .A1(n17382), .A2(img[1482]), .B1(n13798), .B2(img[1354]), 
        .O(n17351) );
  AOI22S U20070 ( .A1(n17864), .A2(img[1994]), .B1(n17383), .B2(img[1866]), 
        .O(n17350) );
  AOI22S U20071 ( .A1(n17347), .A2(img[1226]), .B1(n13787), .B2(img[1098]), 
        .O(n17349) );
  AOI22S U20072 ( .A1(n19036), .A2(img[1738]), .B1(n18201), .B2(img[1610]), 
        .O(n17348) );
  AN4S U20073 ( .I1(n17351), .I2(n17350), .I3(n17349), .I4(n17348), .O(n17352)
         );
  AOI22S U20074 ( .A1(n15506), .A2(img[466]), .B1(n13879), .B2(img[338]), .O(
        n17358) );
  AOI22S U20075 ( .A1(n13788), .A2(img[978]), .B1(n13892), .B2(img[850]), .O(
        n17357) );
  AOI22S U20076 ( .A1(n17354), .A2(img[210]), .B1(n17376), .B2(img[82]), .O(
        n17356) );
  AOI22S U20077 ( .A1(n19641), .A2(img[722]), .B1(n13837), .B2(img[594]), .O(
        n17355) );
  AN4S U20078 ( .I1(n17358), .I2(n17357), .I3(n17356), .I4(n17355), .O(n17365)
         );
  AOI22S U20079 ( .A1(n20109), .A2(img[1490]), .B1(n13798), .B2(img[1362]), 
        .O(n17363) );
  AOI22S U20080 ( .A1(n13801), .A2(img[2002]), .B1(n17383), .B2(img[1874]), 
        .O(n17362) );
  AOI22S U20081 ( .A1(n17359), .A2(img[1234]), .B1(n13787), .B2(img[1106]), 
        .O(n17361) );
  AOI22S U20082 ( .A1(n19023), .A2(img[1746]), .B1(n18201), .B2(img[1618]), 
        .O(n17360) );
  AN4S U20083 ( .I1(n17363), .I2(n17362), .I3(n17361), .I4(n17360), .O(n17364)
         );
  ND2P U20084 ( .I1(n17365), .I2(n17364), .O(n20469) );
  AOI22S U20085 ( .A1(n20476), .A2(n13791), .B1(n13835), .B2(n20469), .O(
        n17366) );
  AN4S U20086 ( .I1(n17369), .I2(n17368), .I3(n17367), .I4(n17366), .O(n17370)
         );
  ND2S U20087 ( .I1(n17371), .I2(n17370), .O(n17432) );
  AOI22S U20088 ( .A1(n20475), .A2(n13839), .B1(n17875), .B2(n20474), .O(
        n17375) );
  AOI22S U20089 ( .A1(n20480), .A2(n20187), .B1(n21062), .B2(n20471), .O(
        n17374) );
  AOI22S U20090 ( .A1(n20489), .A2(n20613), .B1(n17762), .B2(n20481), .O(
        n17373) );
  AOI22S U20091 ( .A1(n20485), .A2(n13830), .B1(n17928), .B2(n20491), .O(
        n17372) );
  AN4S U20092 ( .I1(n17375), .I2(n17374), .I3(n17373), .I4(n17372), .O(n17395)
         );
  AOI22S U20093 ( .A1(n20476), .A2(n20263), .B1(n13847), .B2(n20490), .O(
        n17393) );
  ND2S U20094 ( .I1(n20468), .I2(n20580), .O(n17392) );
  AOI22S U20095 ( .A1(n20102), .A2(img[498]), .B1(n13855), .B2(img[370]), .O(
        n17381) );
  AOI22S U20096 ( .A1(n16515), .A2(img[1010]), .B1(n13880), .B2(img[882]), .O(
        n17380) );
  AOI22S U20097 ( .A1(n17377), .A2(img[242]), .B1(n17376), .B2(img[114]), .O(
        n17379) );
  AOI22S U20098 ( .A1(n19641), .A2(img[754]), .B1(n13898), .B2(img[626]), .O(
        n17378) );
  AOI22S U20099 ( .A1(n17382), .A2(img[1522]), .B1(n17862), .B2(img[1394]), 
        .O(n17387) );
  AOI22S U20100 ( .A1(n17335), .A2(img[2034]), .B1(n17383), .B2(img[1906]), 
        .O(n17386) );
  AOI22S U20101 ( .A1(n13853), .A2(img[1266]), .B1(n18922), .B2(img[1138]), 
        .O(n17385) );
  AOI22S U20102 ( .A1(n19023), .A2(img[1778]), .B1(n18201), .B2(img[1650]), 
        .O(n17384) );
  AN4S U20103 ( .I1(n17387), .I2(n17386), .I3(n17385), .I4(n17384), .O(n17388)
         );
  AOI22S U20104 ( .A1(n20477), .A2(n13804), .B1(n13846), .B2(n20484), .O(
        n17391) );
  AOI22S U20105 ( .A1(n20492), .A2(n19914), .B1(n17938), .B2(n20469), .O(
        n17390) );
  AN4S U20106 ( .I1(n17393), .I2(n17392), .I3(n17391), .I4(n17390), .O(n17394)
         );
  ND2P U20107 ( .I1(n17395), .I2(n17394), .O(n17439) );
  AOI22S U20108 ( .A1(n17432), .A2(n20364), .B1(n20223), .B2(n17439), .O(
        n17435) );
  AOI22S U20109 ( .A1(n19818), .A2(n20484), .B1(n20484), .B2(n22923), .O(
        n17430) );
  NR2 U20110 ( .I1(n17402), .I2(n17401), .O(n17410) );
  AOI22S U20111 ( .A1(n17404), .A2(n13830), .B1(n13839), .B2(n17403), .O(
        n17409) );
  AOI22S U20112 ( .A1(n17407), .A2(n20439), .B1(n17875), .B2(n17406), .O(
        n17408) );
  ND3S U20113 ( .I1(n17410), .I2(n17409), .I3(n17408), .O(n17428) );
  NR2 U20114 ( .I1(n17416), .I2(n17415), .O(n17426) );
  INV1S U20115 ( .I(n17417), .O(n17420) );
  AOI22S U20116 ( .A1(n17420), .A2(n20620), .B1(n13793), .B2(n17419), .O(
        n17425) );
  INV1S U20117 ( .I(n17421), .O(n17423) );
  AOI22S U20118 ( .A1(n17423), .A2(n18040), .B1(n17762), .B2(n17422), .O(
        n17424) );
  ND3 U20119 ( .I1(n17426), .I2(n17425), .I3(n17424), .O(n17427) );
  NR2P U20120 ( .I1(n17428), .I2(n17427), .O(n20388) );
  INV2 U20121 ( .I(n20388), .O(n20358) );
  AOI22S U20122 ( .A1(n20252), .A2(n21225), .B1(n17686), .B2(n20358), .O(
        n17429) );
  AOI12HS U20123 ( .B1(n17432), .B2(n19533), .A1(n17431), .O(n17434) );
  ND2S U20124 ( .I1(n17439), .I2(n20062), .O(n17433) );
  ND2T U20125 ( .I1(n22058), .I2(n20809), .O(n21399) );
  AOI22S U20126 ( .A1(n17439), .A2(n20364), .B1(n19533), .B2(n17439), .O(
        n17442) );
  AOI22S U20127 ( .A1(n19603), .A2(n21225), .B1(n20470), .B2(n22923), .O(
        n17437) );
  ND2S U20128 ( .I1(n20470), .I2(n19818), .O(n17436) );
  ND2S U20129 ( .I1(n17437), .I2(n17436), .O(n17438) );
  AOI12HS U20130 ( .B1(n17439), .B2(n20371), .A1(n17438), .O(n17441) );
  ND2S U20131 ( .I1(n17439), .I2(n19608), .O(n17440) );
  ND3P U20132 ( .I1(n17442), .I2(n17441), .I3(n17440), .O(n21812) );
  AN2P U20133 ( .I1(n21812), .I2(n20809), .O(n20644) );
  ND2S U20134 ( .I1(n17443), .I2(n20644), .O(n17696) );
  AOI22S U20135 ( .A1(n13825), .A2(img[507]), .B1(n13858), .B2(img[379]), .O(
        n17447) );
  AOI22S U20136 ( .A1(n17880), .A2(img[251]), .B1(n19642), .B2(img[123]), .O(
        n17446) );
  AOI22S U20137 ( .A1(n18946), .A2(img[1019]), .B1(n16048), .B2(img[891]), .O(
        n17445) );
  AOI22S U20138 ( .A1(n13886), .A2(img[763]), .B1(n13837), .B2(img[635]), .O(
        n17444) );
  AN4S U20139 ( .I1(n17447), .I2(n17446), .I3(n17445), .I4(n17444), .O(n17453)
         );
  AOI22S U20140 ( .A1(n18729), .A2(img[1275]), .B1(n17885), .B2(img[1147]), 
        .O(n17451) );
  AOI22S U20141 ( .A1(n13786), .A2(img[1787]), .B1(n13796), .B2(img[1659]), 
        .O(n17450) );
  AOI22S U20142 ( .A1(n13823), .A2(img[1531]), .B1(n17862), .B2(img[1403]), 
        .O(n17449) );
  AOI22S U20143 ( .A1(n19411), .A2(img[2043]), .B1(n22928), .B2(img[1915]), 
        .O(n17448) );
  AOI22S U20144 ( .A1(n19603), .A2(n17454), .B1(n19634), .B2(n22923), .O(
        n17456) );
  ND2S U20145 ( .I1(n19634), .I2(n19818), .O(n17455) );
  AOI22S U20146 ( .A1(n15657), .A2(img[491]), .B1(n19709), .B2(img[363]), .O(
        n17460) );
  AOI22S U20147 ( .A1(n14505), .A2(img[1003]), .B1(n13893), .B2(img[875]), .O(
        n17459) );
  AOI22S U20148 ( .A1(n17589), .A2(img[235]), .B1(n17611), .B2(img[107]), .O(
        n17458) );
  AOI22S U20149 ( .A1(n19326), .A2(img[747]), .B1(n13898), .B2(img[619]), .O(
        n17457) );
  AN4S U20150 ( .I1(n17460), .I2(n17459), .I3(n17458), .I4(n17457), .O(n17466)
         );
  AOI22S U20151 ( .A1(n13874), .A2(img[1515]), .B1(n14739), .B2(img[1387]), 
        .O(n17464) );
  BUF1 U20152 ( .I(n22928), .O(n17514) );
  AOI22S U20153 ( .A1(n18958), .A2(img[2027]), .B1(n17617), .B2(img[1899]), 
        .O(n17463) );
  AOI22S U20154 ( .A1(n13783), .A2(img[1259]), .B1(n18623), .B2(img[1131]), 
        .O(n17462) );
  AOI22S U20155 ( .A1(n19036), .A2(img[1771]), .B1(n13796), .B2(img[1643]), 
        .O(n17461) );
  AOI22S U20156 ( .A1(n19343), .A2(img[427]), .B1(n19709), .B2(img[299]), .O(
        n17471) );
  AOI22S U20157 ( .A1(n19037), .A2(img[939]), .B1(n13893), .B2(img[811]), .O(
        n17470) );
  BUF1S U20158 ( .I(n13800), .O(n17467) );
  AOI22S U20159 ( .A1(n17467), .A2(img[171]), .B1(n17611), .B2(img[43]), .O(
        n17469) );
  AOI22S U20160 ( .A1(n13875), .A2(img[683]), .B1(n13837), .B2(img[555]), .O(
        n17468) );
  AN4S U20161 ( .I1(n17471), .I2(n17470), .I3(n17469), .I4(n17468), .O(n17477)
         );
  AOI22S U20162 ( .A1(n17382), .A2(img[1451]), .B1(n17862), .B2(img[1323]), 
        .O(n17475) );
  AOI22S U20163 ( .A1(n14909), .A2(img[1963]), .B1(n17617), .B2(img[1835]), 
        .O(n17474) );
  AOI22S U20164 ( .A1(n13783), .A2(img[1195]), .B1(n13787), .B2(img[1067]), 
        .O(n17473) );
  AOI22S U20165 ( .A1(n19036), .A2(img[1707]), .B1(n13794), .B2(img[1579]), 
        .O(n17472) );
  ND2P U20166 ( .I1(n17477), .I2(n17476), .O(n20413) );
  AOI22S U20167 ( .A1(n20412), .A2(n13839), .B1(n17875), .B2(n20413), .O(
        n17545) );
  AOI22S U20168 ( .A1(n13785), .A2(img[435]), .B1(n13879), .B2(img[307]), .O(
        n17481) );
  AOI22S U20169 ( .A1(n16037), .A2(img[947]), .B1(n13893), .B2(img[819]), .O(
        n17480) );
  BUF1 U20170 ( .I(n13800), .O(n17534) );
  AOI22S U20171 ( .A1(n17534), .A2(img[179]), .B1(n17611), .B2(img[51]), .O(
        n17479) );
  AOI22S U20172 ( .A1(n19326), .A2(img[691]), .B1(n13837), .B2(img[563]), .O(
        n17478) );
  AN4S U20173 ( .I1(n17481), .I2(n17480), .I3(n17479), .I4(n17478), .O(n17487)
         );
  AOI22S U20174 ( .A1(n19193), .A2(img[1459]), .B1(n13845), .B2(img[1331]), 
        .O(n17485) );
  AOI22S U20175 ( .A1(n18773), .A2(img[1971]), .B1(n17617), .B2(img[1843]), 
        .O(n17484) );
  AOI22S U20176 ( .A1(n13783), .A2(img[1203]), .B1(n15800), .B2(img[1075]), 
        .O(n17483) );
  AOI22S U20177 ( .A1(n13870), .A2(img[1715]), .B1(n13832), .B2(img[1587]), 
        .O(n17482) );
  AOI22S U20178 ( .A1(n13785), .A2(img[483]), .B1(n13859), .B2(img[355]), .O(
        n17492) );
  AOI22S U20179 ( .A1(n14189), .A2(img[995]), .B1(n13892), .B2(img[867]), .O(
        n17491) );
  BUF1S U20180 ( .I(n13800), .O(n17488) );
  AOI22S U20181 ( .A1(n17488), .A2(img[227]), .B1(n17611), .B2(img[99]), .O(
        n17490) );
  AOI22S U20182 ( .A1(n19326), .A2(img[739]), .B1(n13797), .B2(img[611]), .O(
        n17489) );
  AOI22S U20183 ( .A1(n19193), .A2(img[1507]), .B1(n13799), .B2(img[1379]), 
        .O(n17496) );
  AOI22S U20184 ( .A1(n13801), .A2(img[2019]), .B1(n17617), .B2(img[1891]), 
        .O(n17495) );
  AOI22S U20185 ( .A1(n13783), .A2(img[1251]), .B1(n17276), .B2(img[1123]), 
        .O(n17494) );
  AOI22S U20186 ( .A1(n13786), .A2(img[1763]), .B1(n13794), .B2(img[1635]), 
        .O(n17493) );
  ND2P U20187 ( .I1(n17498), .I2(n17497), .O(n20411) );
  AOI22S U20188 ( .A1(n20422), .A2(n20187), .B1(n21062), .B2(n20411), .O(
        n17631) );
  AOI22S U20189 ( .A1(n20102), .A2(img[419]), .B1(n13896), .B2(img[291]), .O(
        n17503) );
  AOI22S U20190 ( .A1(n13788), .A2(img[931]), .B1(n13877), .B2(img[803]), .O(
        n17502) );
  BUF1S U20191 ( .I(n13800), .O(n17499) );
  AOI22S U20192 ( .A1(n17499), .A2(img[163]), .B1(n17611), .B2(img[35]), .O(
        n17501) );
  AOI22S U20193 ( .A1(n13875), .A2(img[675]), .B1(n13837), .B2(img[547]), .O(
        n17500) );
  AN4S U20194 ( .I1(n17503), .I2(n17502), .I3(n17501), .I4(n17500), .O(n17509)
         );
  AOI22S U20195 ( .A1(n19193), .A2(img[1443]), .B1(n19182), .B2(img[1315]), 
        .O(n17507) );
  AOI22S U20196 ( .A1(n18958), .A2(img[1955]), .B1(n17617), .B2(img[1827]), 
        .O(n17506) );
  AOI22S U20197 ( .A1(n19856), .A2(img[1187]), .B1(n13787), .B2(img[1059]), 
        .O(n17505) );
  AOI22S U20198 ( .A1(n19036), .A2(img[1699]), .B1(n13794), .B2(img[1571]), 
        .O(n17504) );
  ND2P U20199 ( .I1(n17509), .I2(n17508), .O(n20427) );
  AOI22S U20200 ( .A1(n13785), .A2(img[403]), .B1(n15799), .B2(img[275]), .O(
        n17513) );
  AOI22S U20201 ( .A1(n16037), .A2(img[915]), .B1(n13890), .B2(img[787]), .O(
        n17512) );
  BUF1 U20202 ( .I(n13800), .O(n17578) );
  AOI22S U20203 ( .A1(n17578), .A2(img[147]), .B1(n17611), .B2(img[19]), .O(
        n17511) );
  AOI22S U20204 ( .A1(n19326), .A2(img[659]), .B1(n13797), .B2(img[531]), .O(
        n17510) );
  AN4S U20205 ( .I1(n17513), .I2(n17512), .I3(n17511), .I4(n17510), .O(n17521)
         );
  AOI22S U20206 ( .A1(n17382), .A2(img[1427]), .B1(n19001), .B2(img[1299]), 
        .O(n17519) );
  AOI22S U20207 ( .A1(n17335), .A2(img[1939]), .B1(n17514), .B2(img[1811]), 
        .O(n17518) );
  AOI22S U20208 ( .A1(n13783), .A2(img[1171]), .B1(n19955), .B2(img[1043]), 
        .O(n17517) );
  AOI22S U20209 ( .A1(n19023), .A2(img[1683]), .B1(n13794), .B2(img[1555]), 
        .O(n17516) );
  AN4S U20210 ( .I1(n17519), .I2(n17518), .I3(n17517), .I4(n17516), .O(n17520)
         );
  AOI22S U20211 ( .A1(n20427), .A2(n20613), .B1(n17762), .B2(n20404), .O(
        n17633) );
  AOI22S U20212 ( .A1(n13785), .A2(img[395]), .B1(n15691), .B2(img[267]), .O(
        n17527) );
  AOI22S U20213 ( .A1(n14189), .A2(img[907]), .B1(n13890), .B2(img[779]), .O(
        n17526) );
  BUF1S U20214 ( .I(n13800), .O(n17523) );
  AOI22S U20215 ( .A1(n17523), .A2(img[139]), .B1(n17611), .B2(img[11]), .O(
        n17525) );
  AOI22S U20216 ( .A1(n13875), .A2(img[651]), .B1(n13898), .B2(img[523]), .O(
        n17524) );
  AOI22S U20217 ( .A1(n19193), .A2(img[1419]), .B1(n19001), .B2(img[1291]), 
        .O(n17531) );
  AOI22S U20218 ( .A1(n13841), .A2(img[1931]), .B1(n17617), .B2(img[1803]), 
        .O(n17530) );
  AOI22S U20219 ( .A1(n13827), .A2(img[1163]), .B1(n13787), .B2(img[1035]), 
        .O(n17529) );
  AOI22S U20220 ( .A1(n19036), .A2(img[1675]), .B1(n13832), .B2(img[1547]), 
        .O(n17528) );
  AOI22S U20221 ( .A1(n20102), .A2(img[443]), .B1(n13879), .B2(img[315]), .O(
        n17538) );
  AOI22S U20222 ( .A1(n13788), .A2(img[955]), .B1(n13893), .B2(img[827]), .O(
        n17537) );
  AOI22S U20223 ( .A1(n17534), .A2(img[187]), .B1(n17611), .B2(img[59]), .O(
        n17536) );
  AOI22S U20224 ( .A1(n19326), .A2(img[699]), .B1(n13837), .B2(img[571]), .O(
        n17535) );
  AOI22S U20225 ( .A1(n17382), .A2(img[1467]), .B1(n19182), .B2(img[1339]), 
        .O(n17542) );
  AOI22S U20226 ( .A1(n13801), .A2(img[1979]), .B1(n17617), .B2(img[1851]), 
        .O(n17541) );
  AOI22S U20227 ( .A1(n13783), .A2(img[1211]), .B1(n19417), .B2(img[1083]), 
        .O(n17540) );
  AOI22S U20228 ( .A1(n15751), .A2(img[1723]), .B1(n13832), .B2(img[1595]), 
        .O(n17539) );
  ND2P U20229 ( .I1(n17544), .I2(n17543), .O(n20418) );
  AOI22S U20230 ( .A1(n20419), .A2(n13830), .B1(n17928), .B2(n20418), .O(
        n17632) );
  AN4S U20231 ( .I1(n17545), .I2(n17631), .I3(n17633), .I4(n17632), .O(n17628)
         );
  AOI22S U20232 ( .A1(n13785), .A2(img[459]), .B1(n19709), .B2(img[331]), .O(
        n17549) );
  AOI22S U20233 ( .A1(n18911), .A2(img[971]), .B1(n15653), .B2(img[843]), .O(
        n17548) );
  AOI22S U20234 ( .A1(n17612), .A2(img[203]), .B1(n17611), .B2(img[75]), .O(
        n17547) );
  AOI22S U20235 ( .A1(n19326), .A2(img[715]), .B1(n13797), .B2(img[587]), .O(
        n17546) );
  AOI22S U20236 ( .A1(n19193), .A2(img[1483]), .B1(n19001), .B2(img[1355]), 
        .O(n17554) );
  AOI22S U20237 ( .A1(n17864), .A2(img[1995]), .B1(n17617), .B2(img[1867]), 
        .O(n17553) );
  AOI22S U20238 ( .A1(n13827), .A2(img[1227]), .B1(n17276), .B2(img[1099]), 
        .O(n17552) );
  AOI22S U20239 ( .A1(n19036), .A2(img[1739]), .B1(n17550), .B2(img[1611]), 
        .O(n17551) );
  ND2P U20240 ( .I1(n17556), .I2(n17555), .O(n20414) );
  AOI22S U20241 ( .A1(n13825), .A2(img[387]), .B1(n13858), .B2(img[259]), .O(
        n17560) );
  AOI22S U20242 ( .A1(n16515), .A2(img[899]), .B1(n13861), .B2(img[771]), .O(
        n17559) );
  AOI22S U20243 ( .A1(n13829), .A2(img[131]), .B1(n17611), .B2(img[3]), .O(
        n17558) );
  AOI22S U20244 ( .A1(n19326), .A2(img[643]), .B1(n13797), .B2(img[515]), .O(
        n17557) );
  AN4S U20245 ( .I1(n17560), .I2(n17559), .I3(n17558), .I4(n17557), .O(n17567)
         );
  AOI22S U20246 ( .A1(n19193), .A2(img[1411]), .B1(n18751), .B2(img[1283]), 
        .O(n17565) );
  AOI22S U20247 ( .A1(n17515), .A2(img[1923]), .B1(n17617), .B2(img[1795]), 
        .O(n17564) );
  AOI22S U20248 ( .A1(n13783), .A2(img[1155]), .B1(n18623), .B2(img[1027]), 
        .O(n17563) );
  AOI22S U20249 ( .A1(n19023), .A2(img[1667]), .B1(n17561), .B2(img[1539]), 
        .O(n17562) );
  AOI22S U20250 ( .A1(n20414), .A2(n20263), .B1(n13847), .B2(n20428), .O(
        n17627) );
  AOI22S U20251 ( .A1(n13785), .A2(img[451]), .B1(n13855), .B2(img[323]), .O(
        n17571) );
  AOI22S U20252 ( .A1(n18148), .A2(img[963]), .B1(n13890), .B2(img[835]), .O(
        n17570) );
  BUF1 U20253 ( .I(n13800), .O(n19949) );
  AOI22S U20254 ( .A1(n19949), .A2(img[195]), .B1(n17611), .B2(img[67]), .O(
        n17569) );
  AOI22S U20255 ( .A1(n13875), .A2(img[707]), .B1(n13797), .B2(img[579]), .O(
        n17568) );
  AN4S U20256 ( .I1(n17571), .I2(n17570), .I3(n17569), .I4(n17568), .O(n17577)
         );
  AOI22S U20257 ( .A1(n13823), .A2(img[1475]), .B1(n17862), .B2(img[1347]), 
        .O(n17575) );
  AOI22S U20258 ( .A1(n18958), .A2(img[1987]), .B1(n17617), .B2(img[1859]), 
        .O(n17574) );
  AOI22S U20259 ( .A1(n13783), .A2(img[1219]), .B1(n18623), .B2(img[1091]), 
        .O(n17573) );
  AOI22S U20260 ( .A1(n13867), .A2(img[1731]), .B1(n13794), .B2(img[1603]), 
        .O(n17572) );
  ND2S U20261 ( .I1(n20403), .I2(n20580), .O(n17626) );
  AOI22S U20262 ( .A1(n13876), .A2(img[411]), .B1(n15799), .B2(img[283]), .O(
        n17582) );
  AOI22S U20263 ( .A1(n18946), .A2(img[923]), .B1(n13893), .B2(img[795]), .O(
        n17581) );
  AOI22S U20264 ( .A1(n17578), .A2(img[155]), .B1(n17611), .B2(img[27]), .O(
        n17580) );
  AOI22S U20265 ( .A1(n19326), .A2(img[667]), .B1(n13837), .B2(img[539]), .O(
        n17579) );
  AN4S U20266 ( .I1(n17582), .I2(n17581), .I3(n17580), .I4(n17579), .O(n17588)
         );
  AOI22S U20267 ( .A1(n19193), .A2(img[1435]), .B1(n13845), .B2(img[1307]), 
        .O(n17586) );
  AOI22S U20268 ( .A1(n18996), .A2(img[1947]), .B1(n17617), .B2(img[1819]), 
        .O(n17585) );
  AOI22S U20269 ( .A1(n18729), .A2(img[1179]), .B1(n13802), .B2(img[1051]), 
        .O(n17584) );
  AOI22S U20270 ( .A1(n13786), .A2(img[1691]), .B1(n13832), .B2(img[1563]), 
        .O(n17583) );
  AN4S U20271 ( .I1(n17586), .I2(n17585), .I3(n17584), .I4(n17583), .O(n17587)
         );
  AOI22S U20272 ( .A1(n13785), .A2(img[499]), .B1(n13855), .B2(img[371]), .O(
        n17593) );
  AOI22S U20273 ( .A1(n18946), .A2(img[1011]), .B1(n13889), .B2(img[883]), .O(
        n17592) );
  AOI22S U20274 ( .A1(n17589), .A2(img[243]), .B1(n17611), .B2(img[115]), .O(
        n17591) );
  AOI22S U20275 ( .A1(n13875), .A2(img[755]), .B1(n13837), .B2(img[627]), .O(
        n17590) );
  AN4 U20276 ( .I1(n17593), .I2(n17592), .I3(n17591), .I4(n17590), .O(n17599)
         );
  AOI22S U20277 ( .A1(n18837), .A2(img[1523]), .B1(n17827), .B2(img[1395]), 
        .O(n17597) );
  AOI22S U20278 ( .A1(n13801), .A2(img[2035]), .B1(n17617), .B2(img[1907]), 
        .O(n17596) );
  AOI22S U20279 ( .A1(n18897), .A2(img[1267]), .B1(n15800), .B2(img[1139]), 
        .O(n17595) );
  AOI22S U20280 ( .A1(n20038), .A2(img[1779]), .B1(n13794), .B2(img[1651]), 
        .O(n17594) );
  ND2P U20281 ( .I1(n17599), .I2(n17598), .O(n19625) );
  AOI22S U20282 ( .A1(n20426), .A2(n13804), .B1(n13846), .B2(n19625), .O(
        n17625) );
  AOI22S U20283 ( .A1(n13785), .A2(img[475]), .B1(n19709), .B2(img[347]), .O(
        n17604) );
  AOI22S U20284 ( .A1(n18911), .A2(img[987]), .B1(n13893), .B2(img[859]), .O(
        n17603) );
  BUF1S U20285 ( .I(n13800), .O(n17600) );
  AOI22S U20286 ( .A1(n17600), .A2(img[219]), .B1(n17611), .B2(img[91]), .O(
        n17602) );
  AOI22S U20287 ( .A1(n13875), .A2(img[731]), .B1(n13797), .B2(img[603]), .O(
        n17601) );
  AOI22S U20288 ( .A1(n15630), .A2(img[1499]), .B1(n17827), .B2(img[1371]), 
        .O(n17608) );
  AOI22S U20289 ( .A1(n18996), .A2(img[2011]), .B1(n17617), .B2(img[1883]), 
        .O(n17607) );
  AOI22S U20290 ( .A1(n19856), .A2(img[1243]), .B1(n19955), .B2(img[1115]), 
        .O(n17606) );
  AOI22S U20291 ( .A1(n13786), .A2(img[1755]), .B1(n13796), .B2(img[1627]), 
        .O(n17605) );
  ND2P U20292 ( .I1(n17610), .I2(n17609), .O(n20429) );
  AOI22S U20293 ( .A1(n20102), .A2(img[467]), .B1(n19709), .B2(img[339]), .O(
        n17616) );
  AOI22S U20294 ( .A1(n13788), .A2(img[979]), .B1(n13880), .B2(img[851]), .O(
        n17615) );
  AOI22S U20295 ( .A1(n17612), .A2(img[211]), .B1(n17611), .B2(img[83]), .O(
        n17614) );
  AOI22S U20296 ( .A1(n19326), .A2(img[723]), .B1(n13797), .B2(img[595]), .O(
        n17613) );
  AOI22S U20297 ( .A1(n19193), .A2(img[1491]), .B1(n13799), .B2(img[1363]), 
        .O(n17621) );
  AOI22S U20298 ( .A1(n17335), .A2(img[2003]), .B1(n17617), .B2(img[1875]), 
        .O(n17620) );
  AOI22S U20299 ( .A1(n17088), .A2(img[1235]), .B1(n19417), .B2(img[1107]), 
        .O(n17619) );
  AOI22S U20300 ( .A1(n19215), .A2(img[1747]), .B1(n13794), .B2(img[1619]), 
        .O(n17618) );
  ND2P U20301 ( .I1(n17623), .I2(n17622), .O(n20407) );
  AOI22S U20302 ( .A1(n20429), .A2(n13835), .B1(n17938), .B2(n20407), .O(
        n17624) );
  AN4S U20303 ( .I1(n17627), .I2(n17626), .I3(n17625), .I4(n17624), .O(n17638)
         );
  AOI22S U20304 ( .A1(n17653), .A2(n19533), .B1(n20314), .B2(n17653), .O(
        n17641) );
  ND2S U20305 ( .I1(n20412), .I2(n13839), .O(n17630) );
  ND2S U20306 ( .I1(n20413), .I2(n17875), .O(n17629) );
  ND3S U20307 ( .I1(n17631), .I2(n17630), .I3(n17629), .O(n17635) );
  ND2S U20308 ( .I1(n17633), .I2(n17632), .O(n17634) );
  NR2 U20309 ( .I1(n17635), .I2(n17634), .O(n17637) );
  AO12 U20310 ( .B1(n17638), .B2(n17637), .A1(n17636), .O(n17642) );
  INV1S U20311 ( .I(n17642), .O(n17639) );
  AOI12HS U20312 ( .B1(n20364), .B2(n17653), .A1(n17639), .O(n17640) );
  ND3HT U20313 ( .I1(n13932), .I2(n17641), .I3(n17640), .O(n21811) );
  AN2T U20314 ( .I1(n21811), .I2(n20809), .O(n20503) );
  OR2 U20315 ( .I1(n13822), .I2(n17642), .O(n17694) );
  AOI22S U20316 ( .A1(n20411), .A2(n13839), .B1(n17875), .B2(n20427), .O(
        n17646) );
  AOI22S U20317 ( .A1(n20429), .A2(n19483), .B1(n20187), .B2(n20413), .O(
        n17645) );
  AOI22S U20318 ( .A1(n20426), .A2(n20613), .B1(n17762), .B2(n20419), .O(
        n17644) );
  AOI22S U20319 ( .A1(n20428), .A2(n13830), .B1(n17928), .B2(n20422), .O(
        n17643) );
  AN4S U20320 ( .I1(n17646), .I2(n17645), .I3(n17644), .I4(n17643), .O(n17652)
         );
  AOI22S U20321 ( .A1(n20403), .A2(n20263), .B1(n13847), .B2(n19634), .O(
        n17650) );
  ND2S U20322 ( .I1(n20418), .I2(n20560), .O(n17649) );
  AOI22S U20323 ( .A1(n20412), .A2(n13846), .B1(n20438), .B2(n20404), .O(
        n17648) );
  AOI22S U20324 ( .A1(n20414), .A2(n13791), .B1(n13835), .B2(n20407), .O(
        n17647) );
  AN4S U20325 ( .I1(n17650), .I2(n17649), .I3(n17648), .I4(n17647), .O(n17651)
         );
  ND2S U20326 ( .I1(n17652), .I2(n17651), .O(n17691) );
  AOI22S U20327 ( .A1(n17653), .A2(n20223), .B1(n20364), .B2(n17691), .O(
        n17693) );
  ND2S U20328 ( .I1(n19625), .I2(n22923), .O(n17689) );
  MOAI1 U20329 ( .A1(n17655), .A2(n15142), .B1(n17654), .B2(n17875), .O(n17661) );
  OAI22S U20330 ( .A1(n17659), .A2(n17658), .B1(n17657), .B2(n17656), .O(
        n17660) );
  AOI22S U20331 ( .A1(n17663), .A2(n19483), .B1(n20438), .B2(n17662), .O(
        n17667) );
  AOI22S U20332 ( .A1(n17665), .A2(n13791), .B1(n17664), .B2(n20263), .O(
        n17666) );
  NR2 U20333 ( .I1(n17674), .I2(n17673), .O(n17683) );
  INV1S U20334 ( .I(n17675), .O(n17676) );
  AOI22S U20335 ( .A1(n13839), .A2(n17677), .B1(n17676), .B2(n20124), .O(
        n17682) );
  MAOI1S U20336 ( .A1(n20969), .A2(n17680), .B1(n13945), .B2(n17678), .O(
        n17681) );
  ND3 U20337 ( .I1(n17683), .I2(n17682), .I3(n17681), .O(n17684) );
  INV2 U20338 ( .I(n20679), .O(n20357) );
  ND2S U20339 ( .I1(n17686), .I2(n20357), .O(n17687) );
  ND3 U20340 ( .I1(n17689), .I2(n17688), .I3(n17687), .O(n17690) );
  AOI12H U20341 ( .B1(n17691), .B2(n19533), .A1(n17690), .O(n17692) );
  ND3HT U20342 ( .I1(n17694), .I2(n17693), .I3(n17692), .O(n22059) );
  OAI112HS U20343 ( .C1(n17697), .C2(n29491), .A1(n17696), .B1(n17695), .O(
        n17962) );
  ND2F U20344 ( .I1(n22059), .I2(n20809), .O(n21403) );
  AOI22S U20345 ( .A1(n19343), .A2(img[492]), .B1(n15799), .B2(img[364]), .O(
        n17701) );
  AOI22S U20346 ( .A1(n18946), .A2(img[1004]), .B1(n13889), .B2(img[876]), .O(
        n17700) );
  AOI22S U20347 ( .A1(n17330), .A2(img[236]), .B1(n17611), .B2(img[108]), .O(
        n17699) );
  AOI22S U20348 ( .A1(n17835), .A2(img[748]), .B1(n13797), .B2(img[620]), .O(
        n17698) );
  AN4S U20349 ( .I1(n17701), .I2(n17700), .I3(n17699), .I4(n17698), .O(n17707)
         );
  AOI22S U20350 ( .A1(n15630), .A2(img[1516]), .B1(n17862), .B2(img[1388]), 
        .O(n17705) );
  AOI22S U20351 ( .A1(n13841), .A2(img[2028]), .B1(n17863), .B2(img[1900]), 
        .O(n17704) );
  AOI22S U20352 ( .A1(n14392), .A2(img[1260]), .B1(n17840), .B2(img[1132]), 
        .O(n17703) );
  AOI22S U20353 ( .A1(n19023), .A2(img[1772]), .B1(n13794), .B2(img[1644]), 
        .O(n17702) );
  AOI22S U20354 ( .A1(n13883), .A2(img[428]), .B1(n19709), .B2(img[300]), .O(
        n17711) );
  AOI22S U20355 ( .A1(n16515), .A2(img[940]), .B1(n16048), .B2(img[812]), .O(
        n17710) );
  AOI22S U20356 ( .A1(n17249), .A2(img[172]), .B1(n17611), .B2(img[44]), .O(
        n17709) );
  AOI22S U20357 ( .A1(n13784), .A2(img[684]), .B1(n13837), .B2(img[556]), .O(
        n17708) );
  AN4S U20358 ( .I1(n17711), .I2(n17710), .I3(n17709), .I4(n17708), .O(n17718)
         );
  AOI22S U20359 ( .A1(n19193), .A2(img[1452]), .B1(n13798), .B2(img[1324]), 
        .O(n17716) );
  AOI22S U20360 ( .A1(n17886), .A2(img[1964]), .B1(n17863), .B2(img[1836]), 
        .O(n17715) );
  AOI22S U20361 ( .A1(n17088), .A2(img[1196]), .B1(n17712), .B2(img[1068]), 
        .O(n17714) );
  AOI22S U20362 ( .A1(n13867), .A2(img[1708]), .B1(n13832), .B2(img[1580]), 
        .O(n17713) );
  AOI22S U20363 ( .A1(n20512), .A2(n13839), .B1(n17875), .B2(n20513), .O(
        n17904) );
  AOI22S U20364 ( .A1(n15506), .A2(img[436]), .B1(n19709), .B2(img[308]), .O(
        n17722) );
  AOI22S U20365 ( .A1(n16515), .A2(img[948]), .B1(n13893), .B2(img[820]), .O(
        n17721) );
  AOI22S U20366 ( .A1(n17197), .A2(img[180]), .B1(n17611), .B2(img[52]), .O(
        n17720) );
  AOI22S U20367 ( .A1(n13875), .A2(img[692]), .B1(n13797), .B2(img[564]), .O(
        n17719) );
  AOI22S U20368 ( .A1(n19193), .A2(img[1460]), .B1(n13798), .B2(img[1332]), 
        .O(n17726) );
  AOI22S U20369 ( .A1(n13803), .A2(img[1972]), .B1(n17863), .B2(img[1844]), 
        .O(n17725) );
  AOI22S U20370 ( .A1(n19856), .A2(img[1204]), .B1(n13802), .B2(img[1076]), 
        .O(n17724) );
  AOI22S U20371 ( .A1(n13863), .A2(img[1716]), .B1(n13796), .B2(img[1588]), 
        .O(n17723) );
  AOI22S U20372 ( .A1(n19343), .A2(img[484]), .B1(n13879), .B2(img[356]), .O(
        n17734) );
  AOI22S U20373 ( .A1(n13788), .A2(img[996]), .B1(n13893), .B2(img[868]), .O(
        n17733) );
  AOI22S U20374 ( .A1(n17729), .A2(img[228]), .B1(n20103), .B2(img[100]), .O(
        n17732) );
  AOI22S U20375 ( .A1(n17730), .A2(img[740]), .B1(n13837), .B2(img[612]), .O(
        n17731) );
  AN4S U20376 ( .I1(n17734), .I2(n17733), .I3(n17732), .I4(n17731), .O(n17740)
         );
  AOI22S U20377 ( .A1(n15630), .A2(img[1508]), .B1(n17862), .B2(img[1380]), 
        .O(n17738) );
  AOI22S U20378 ( .A1(n17886), .A2(img[2020]), .B1(n17863), .B2(img[1892]), 
        .O(n17737) );
  AOI22S U20379 ( .A1(n13853), .A2(img[1252]), .B1(n13802), .B2(img[1124]), 
        .O(n17736) );
  AOI22S U20380 ( .A1(n19023), .A2(img[1764]), .B1(n13794), .B2(img[1636]), 
        .O(n17735) );
  AOI22S U20381 ( .A1(n20526), .A2(n20963), .B1(n21062), .B2(n20511), .O(
        n17903) );
  AOI22S U20382 ( .A1(n13785), .A2(img[420]), .B1(n13879), .B2(img[292]), .O(
        n17744) );
  AOI22S U20383 ( .A1(n16515), .A2(img[932]), .B1(n13890), .B2(img[804]), .O(
        n17743) );
  AOI22S U20384 ( .A1(n17218), .A2(img[164]), .B1(n17611), .B2(img[36]), .O(
        n17742) );
  AOI22S U20385 ( .A1(n19641), .A2(img[676]), .B1(n13797), .B2(img[548]), .O(
        n17741) );
  AN4S U20386 ( .I1(n17744), .I2(n17743), .I3(n17742), .I4(n17741), .O(n17751)
         );
  AOI22S U20387 ( .A1(n19193), .A2(img[1444]), .B1(n13798), .B2(img[1316]), 
        .O(n17749) );
  AOI22S U20388 ( .A1(n17816), .A2(img[1956]), .B1(n17863), .B2(img[1828]), 
        .O(n17748) );
  AOI22S U20389 ( .A1(n17254), .A2(img[1188]), .B1(n17745), .B2(img[1060]), 
        .O(n17747) );
  AOI22S U20390 ( .A1(n19215), .A2(img[1700]), .B1(n13794), .B2(img[1572]), 
        .O(n17746) );
  ND2P U20391 ( .I1(n17751), .I2(n17750), .O(n20519) );
  AOI22S U20392 ( .A1(n13825), .A2(img[404]), .B1(n13896), .B2(img[276]), .O(
        n17755) );
  AOI22S U20393 ( .A1(n18911), .A2(img[916]), .B1(n13893), .B2(img[788]), .O(
        n17754) );
  AOI22S U20394 ( .A1(n19266), .A2(img[148]), .B1(n17611), .B2(img[20]), .O(
        n17753) );
  AOI22S U20395 ( .A1(n13784), .A2(img[660]), .B1(n13837), .B2(img[532]), .O(
        n17752) );
  AN4S U20396 ( .I1(n17755), .I2(n17754), .I3(n17753), .I4(n17752), .O(n17761)
         );
  AOI22S U20397 ( .A1(n19193), .A2(img[1428]), .B1(n17827), .B2(img[1300]), 
        .O(n17759) );
  AOI22S U20398 ( .A1(n17816), .A2(img[1940]), .B1(n17863), .B2(img[1812]), 
        .O(n17758) );
  AOI22S U20399 ( .A1(n13853), .A2(img[1172]), .B1(n18922), .B2(img[1044]), 
        .O(n17757) );
  AOI22S U20400 ( .A1(n19215), .A2(img[1684]), .B1(n17561), .B2(img[1556]), 
        .O(n17756) );
  AN4S U20401 ( .I1(n17759), .I2(n17758), .I3(n17757), .I4(n17756), .O(n17760)
         );
  AOI22S U20402 ( .A1(n20519), .A2(n20613), .B1(n17762), .B2(n20507), .O(
        n17787) );
  AOI22S U20403 ( .A1(n13876), .A2(img[396]), .B1(n15799), .B2(img[268]), .O(
        n17766) );
  AOI22S U20404 ( .A1(n13788), .A2(img[908]), .B1(n13861), .B2(img[780]), .O(
        n17765) );
  AOI22S U20405 ( .A1(n13800), .A2(img[140]), .B1(n17376), .B2(img[12]), .O(
        n17764) );
  AOI22S U20406 ( .A1(n19252), .A2(img[652]), .B1(n13837), .B2(img[524]), .O(
        n17763) );
  AN4S U20407 ( .I1(n17766), .I2(n17765), .I3(n17764), .I4(n17763), .O(n17773)
         );
  AOI22S U20408 ( .A1(n15630), .A2(img[1420]), .B1(n13798), .B2(img[1292]), 
        .O(n17771) );
  AOI22S U20409 ( .A1(n19411), .A2(img[1932]), .B1(n17863), .B2(img[1804]), 
        .O(n17770) );
  AOI22S U20410 ( .A1(n16635), .A2(img[1164]), .B1(n17767), .B2(img[1036]), 
        .O(n17769) );
  AOI22S U20411 ( .A1(n19036), .A2(img[1676]), .B1(n18201), .B2(img[1548]), 
        .O(n17768) );
  ND2P U20412 ( .I1(n17773), .I2(n17772), .O(n20525) );
  AOI22S U20413 ( .A1(n15506), .A2(img[444]), .B1(n13855), .B2(img[316]), .O(
        n17777) );
  AOI22S U20414 ( .A1(n20110), .A2(img[956]), .B1(n13889), .B2(img[828]), .O(
        n17776) );
  AOI22S U20415 ( .A1(n17612), .A2(img[188]), .B1(n13836), .B2(img[60]), .O(
        n17775) );
  AOI22S U20416 ( .A1(n13875), .A2(img[700]), .B1(n13837), .B2(img[572]), .O(
        n17774) );
  AN4S U20417 ( .I1(n17777), .I2(n17776), .I3(n17775), .I4(n17774), .O(n17785)
         );
  AOI22S U20418 ( .A1(n19411), .A2(img[1980]), .B1(n17863), .B2(img[1852]), 
        .O(n17782) );
  AOI22S U20419 ( .A1(n13783), .A2(img[1212]), .B1(n13802), .B2(img[1084]), 
        .O(n17781) );
  AOI22S U20420 ( .A1(n13867), .A2(img[1724]), .B1(n13794), .B2(img[1596]), 
        .O(n17780) );
  AN4S U20421 ( .I1(n17783), .I2(n17782), .I3(n17781), .I4(n17780), .O(n17784)
         );
  AOI22S U20422 ( .A1(n20525), .A2(n13830), .B1(n17928), .B2(n20523), .O(
        n17786) );
  AN4S U20423 ( .I1(n17904), .I2(n17903), .I3(n17787), .I4(n17786), .O(n17874)
         );
  AOI22S U20424 ( .A1(n18681), .A2(img[460]), .B1(n13859), .B2(img[332]), .O(
        n17792) );
  AOI22S U20425 ( .A1(n18946), .A2(img[972]), .B1(n16048), .B2(img[844]), .O(
        n17791) );
  AOI22S U20426 ( .A1(n17788), .A2(img[204]), .B1(n19388), .B2(img[76]), .O(
        n17790) );
  AOI22S U20427 ( .A1(n16348), .A2(img[716]), .B1(n13797), .B2(img[588]), .O(
        n17789) );
  AN4S U20428 ( .I1(n17792), .I2(n17791), .I3(n17790), .I4(n17789), .O(n17799)
         );
  AOI22S U20429 ( .A1(n19193), .A2(img[1484]), .B1(n17862), .B2(img[1356]), 
        .O(n17797) );
  AOI22S U20430 ( .A1(n18996), .A2(img[1996]), .B1(n17863), .B2(img[1868]), 
        .O(n17796) );
  AOI22S U20431 ( .A1(n15315), .A2(img[1228]), .B1(n20198), .B2(img[1100]), 
        .O(n17795) );
  AOI22S U20432 ( .A1(n19036), .A2(img[1740]), .B1(n13794), .B2(img[1612]), 
        .O(n17794) );
  AOI22S U20433 ( .A1(n20032), .A2(img[388]), .B1(n13896), .B2(img[260]), .O(
        n17803) );
  AOI22S U20434 ( .A1(n18946), .A2(img[900]), .B1(n15653), .B2(img[772]), .O(
        n17802) );
  AOI22S U20435 ( .A1(n17249), .A2(img[132]), .B1(n20103), .B2(img[4]), .O(
        n17801) );
  AOI22S U20436 ( .A1(n19641), .A2(img[644]), .B1(n13898), .B2(img[516]), .O(
        n17800) );
  AN4S U20437 ( .I1(n17803), .I2(n17802), .I3(n17801), .I4(n17800), .O(n17809)
         );
  AOI22S U20438 ( .A1(n19193), .A2(img[1412]), .B1(n17827), .B2(img[1284]), 
        .O(n17807) );
  AOI22S U20439 ( .A1(n20104), .A2(img[1924]), .B1(n17863), .B2(img[1796]), 
        .O(n17806) );
  AOI22S U20440 ( .A1(n13824), .A2(img[1156]), .B1(n18838), .B2(img[1028]), 
        .O(n17805) );
  AOI22S U20441 ( .A1(n19023), .A2(img[1668]), .B1(n13796), .B2(img[1540]), 
        .O(n17804) );
  AOI22S U20442 ( .A1(n20514), .A2(n20263), .B1(n13847), .B2(n20521), .O(
        n17872) );
  AOI22S U20443 ( .A1(n13785), .A2(img[452]), .B1(n13859), .B2(img[324]), .O(
        n17815) );
  AOI22S U20444 ( .A1(n16515), .A2(img[964]), .B1(n13861), .B2(img[836]), .O(
        n17814) );
  AOI22S U20445 ( .A1(n17811), .A2(img[196]), .B1(n20103), .B2(img[68]), .O(
        n17813) );
  AOI22S U20446 ( .A1(n19641), .A2(img[708]), .B1(n13837), .B2(img[580]), .O(
        n17812) );
  AN4S U20447 ( .I1(n17815), .I2(n17814), .I3(n17813), .I4(n17812), .O(n17822)
         );
  AOI22S U20448 ( .A1(n19193), .A2(img[1476]), .B1(n13798), .B2(img[1348]), 
        .O(n17820) );
  AOI22S U20449 ( .A1(n14909), .A2(img[1988]), .B1(n17863), .B2(img[1860]), 
        .O(n17819) );
  AOI22S U20450 ( .A1(n13783), .A2(img[1220]), .B1(n13792), .B2(img[1092]), 
        .O(n17818) );
  AOI22S U20451 ( .A1(n19036), .A2(img[1732]), .B1(n13794), .B2(img[1604]), 
        .O(n17817) );
  AN4S U20452 ( .I1(n17820), .I2(n17819), .I3(n17818), .I4(n17817), .O(n17821)
         );
  ND2S U20453 ( .I1(n20508), .I2(n20524), .O(n17908) );
  AOI22S U20454 ( .A1(n13785), .A2(img[412]), .B1(n13896), .B2(img[284]), .O(
        n17826) );
  AOI22S U20455 ( .A1(n13788), .A2(img[924]), .B1(n13889), .B2(img[796]), .O(
        n17825) );
  AOI22S U20456 ( .A1(n17330), .A2(img[156]), .B1(n17611), .B2(img[28]), .O(
        n17824) );
  AOI22S U20457 ( .A1(n13784), .A2(img[668]), .B1(n13837), .B2(img[540]), .O(
        n17823) );
  AN4S U20458 ( .I1(n17826), .I2(n17825), .I3(n17824), .I4(n17823), .O(n17834)
         );
  AOI22S U20459 ( .A1(n19193), .A2(img[1436]), .B1(n17827), .B2(img[1308]), 
        .O(n17832) );
  AOI22S U20460 ( .A1(n18983), .A2(img[1948]), .B1(n17863), .B2(img[1820]), 
        .O(n17831) );
  AOI22S U20461 ( .A1(n13853), .A2(img[1180]), .B1(n18922), .B2(img[1052]), 
        .O(n17830) );
  AOI22S U20462 ( .A1(n19036), .A2(img[1692]), .B1(n18201), .B2(img[1564]), 
        .O(n17829) );
  AOI22S U20463 ( .A1(n19343), .A2(img[500]), .B1(n13896), .B2(img[372]), .O(
        n17839) );
  AOI22S U20464 ( .A1(n18911), .A2(img[1012]), .B1(n13889), .B2(img[884]), .O(
        n17838) );
  AOI22S U20465 ( .A1(n17197), .A2(img[244]), .B1(n17611), .B2(img[116]), .O(
        n17837) );
  AOI22S U20466 ( .A1(n17835), .A2(img[756]), .B1(n13797), .B2(img[628]), .O(
        n17836) );
  AN4S U20467 ( .I1(n17839), .I2(n17838), .I3(n17837), .I4(n17836), .O(n17846)
         );
  AOI22S U20468 ( .A1(n15630), .A2(img[1524]), .B1(n17862), .B2(img[1396]), 
        .O(n17844) );
  AOI22S U20469 ( .A1(n17886), .A2(img[2036]), .B1(n17863), .B2(img[1908]), 
        .O(n17843) );
  AOI22S U20470 ( .A1(n15315), .A2(img[1268]), .B1(n17840), .B2(img[1140]), 
        .O(n17842) );
  AOI22S U20471 ( .A1(n19036), .A2(img[1780]), .B1(n13794), .B2(img[1652]), 
        .O(n17841) );
  AOI22S U20472 ( .A1(n20520), .A2(n13804), .B1(n13846), .B2(n20527), .O(
        n17911) );
  AOI22S U20473 ( .A1(n13785), .A2(img[476]), .B1(n13858), .B2(img[348]), .O(
        n17850) );
  AOI22S U20474 ( .A1(n14189), .A2(img[988]), .B1(n16048), .B2(img[860]), .O(
        n17849) );
  AOI22S U20475 ( .A1(n17857), .A2(img[220]), .B1(n17611), .B2(img[92]), .O(
        n17848) );
  AOI22S U20476 ( .A1(n19641), .A2(img[732]), .B1(n13837), .B2(img[604]), .O(
        n17847) );
  AN4S U20477 ( .I1(n17850), .I2(n17849), .I3(n17848), .I4(n17847), .O(n17856)
         );
  AOI22S U20478 ( .A1(n13823), .A2(img[1500]), .B1(n17862), .B2(img[1372]), 
        .O(n17854) );
  AOI22S U20479 ( .A1(n18983), .A2(img[2012]), .B1(n17863), .B2(img[1884]), 
        .O(n17853) );
  AOI22S U20480 ( .A1(n17312), .A2(img[1244]), .B1(n17865), .B2(img[1116]), 
        .O(n17852) );
  AOI22S U20481 ( .A1(n19036), .A2(img[1756]), .B1(n13794), .B2(img[1628]), 
        .O(n17851) );
  AN4 U20482 ( .I1(n17854), .I2(n17853), .I3(n17852), .I4(n17851), .O(n17855)
         );
  AOI22S U20483 ( .A1(n15657), .A2(img[468]), .B1(n19709), .B2(img[340]), .O(
        n17861) );
  AOI22S U20484 ( .A1(n18935), .A2(img[980]), .B1(n13877), .B2(img[852]), .O(
        n17860) );
  AOI22S U20485 ( .A1(n17857), .A2(img[212]), .B1(n17376), .B2(img[84]), .O(
        n17859) );
  AOI22S U20486 ( .A1(n19641), .A2(img[724]), .B1(n13837), .B2(img[596]), .O(
        n17858) );
  AN4S U20487 ( .I1(n17861), .I2(n17860), .I3(n17859), .I4(n17858), .O(n17871)
         );
  AOI22S U20488 ( .A1(n19193), .A2(img[1492]), .B1(n17862), .B2(img[1364]), 
        .O(n17869) );
  AOI22S U20489 ( .A1(n13833), .A2(img[2004]), .B1(n17863), .B2(img[1876]), 
        .O(n17868) );
  AOI22S U20490 ( .A1(n13783), .A2(img[1236]), .B1(n17865), .B2(img[1108]), 
        .O(n17867) );
  AOI22S U20491 ( .A1(n19036), .A2(img[1748]), .B1(n17561), .B2(img[1620]), 
        .O(n17866) );
  AN4S U20492 ( .I1(n17869), .I2(n17868), .I3(n17867), .I4(n17866), .O(n17870)
         );
  AOI22S U20493 ( .A1(n20522), .A2(n13835), .B1(n17938), .B2(n20510), .O(
        n17910) );
  ND2 U20494 ( .I1(n17874), .I2(n17873), .O(n17957) );
  AOI22S U20495 ( .A1(n20511), .A2(n13839), .B1(n17875), .B2(n20519), .O(
        n17879) );
  AOI22S U20496 ( .A1(n20522), .A2(n19483), .B1(n20187), .B2(n20513), .O(
        n17878) );
  AOI22S U20497 ( .A1(n20520), .A2(n20613), .B1(n17762), .B2(n20525), .O(
        n17877) );
  AOI22S U20498 ( .A1(n20521), .A2(n13830), .B1(n17928), .B2(n20526), .O(
        n17876) );
  AN4S U20499 ( .I1(n17879), .I2(n17878), .I3(n17877), .I4(n17876), .O(n17898)
         );
  AOI22S U20500 ( .A1(n13825), .A2(img[508]), .B1(n13858), .B2(img[380]), .O(
        n17884) );
  AOI22S U20501 ( .A1(n17880), .A2(img[252]), .B1(n19642), .B2(img[124]), .O(
        n17883) );
  AOI22S U20502 ( .A1(n18946), .A2(img[1020]), .B1(n13889), .B2(img[892]), .O(
        n17882) );
  AOI22S U20503 ( .A1(n13886), .A2(img[764]), .B1(n13837), .B2(img[636]), .O(
        n17881) );
  AN4S U20504 ( .I1(n17884), .I2(n17883), .I3(n17882), .I4(n17881), .O(n17892)
         );
  AOI22S U20505 ( .A1(n18923), .A2(img[1276]), .B1(n17885), .B2(img[1148]), 
        .O(n17890) );
  AOI22S U20506 ( .A1(n19215), .A2(img[1788]), .B1(n13794), .B2(img[1660]), 
        .O(n17889) );
  AOI22S U20507 ( .A1(n17382), .A2(img[1532]), .B1(n13845), .B2(img[1404]), 
        .O(n17888) );
  AOI22S U20508 ( .A1(n17515), .A2(img[2044]), .B1(n22928), .B2(img[1916]), 
        .O(n17887) );
  AN4S U20509 ( .I1(n17890), .I2(n17889), .I3(n17888), .I4(n17887), .O(n17891)
         );
  AOI22S U20510 ( .A1(n20508), .A2(n20439), .B1(n13847), .B2(n20509), .O(
        n17896) );
  ND2S U20511 ( .I1(n20523), .I2(n20580), .O(n17895) );
  AOI22S U20512 ( .A1(n20512), .A2(n13846), .B1(n20438), .B2(n20507), .O(
        n17894) );
  AOI22S U20513 ( .A1(n20514), .A2(n13791), .B1(n13835), .B2(n20510), .O(
        n17893) );
  AN4S U20514 ( .I1(n17896), .I2(n17895), .I3(n17894), .I4(n17893), .O(n17897)
         );
  ND2S U20515 ( .I1(n17898), .I2(n17897), .O(n17949) );
  AOI22S U20516 ( .A1(n17957), .A2(n20223), .B1(n20364), .B2(n17949), .O(
        n17952) );
  ND2S U20517 ( .I1(n20519), .I2(n20613), .O(n17902) );
  ND2S U20518 ( .I1(n20507), .I2(n17762), .O(n17901) );
  ND2S U20519 ( .I1(n20525), .I2(n13830), .O(n17900) );
  ND2S U20520 ( .I1(n20523), .I2(n17928), .O(n17899) );
  AN4S U20521 ( .I1(n17902), .I2(n17901), .I3(n17900), .I4(n17899), .O(n17905)
         );
  ND3S U20522 ( .I1(n17905), .I2(n17904), .I3(n17903), .O(n17914) );
  ND2S U20523 ( .I1(n20514), .I2(n20263), .O(n17907) );
  ND2S U20524 ( .I1(n20521), .I2(n13847), .O(n17906) );
  ND3S U20525 ( .I1(n17908), .I2(n17907), .I3(n17906), .O(n17909) );
  INV1S U20526 ( .I(n17909), .O(n17912) );
  ND3S U20527 ( .I1(n17912), .I2(n17911), .I3(n17910), .O(n17913) );
  OAI12HS U20528 ( .B1(n17914), .B2(n17913), .A1(n19608), .O(n17958) );
  OR2 U20529 ( .I1(n13822), .I2(n17958), .O(n17951) );
  ND2S U20530 ( .I1(n20527), .I2(n22923), .O(n17947) );
  MOAI1 U20531 ( .A1(n17918), .A2(n15142), .B1(n17917), .B2(n17762), .O(n17926) );
  AOI22S U20532 ( .A1(n17920), .A2(n17875), .B1(n20124), .B2(n17919), .O(
        n17923) );
  ND2S U20533 ( .I1(n17921), .I2(n20969), .O(n17922) );
  OAI112HS U20534 ( .C1(n17924), .C2(n13929), .A1(n17923), .B1(n17922), .O(
        n17925) );
  NR2 U20535 ( .I1(n17935), .I2(n17934), .O(n17944) );
  MOAI1 U20536 ( .A1(n17940), .A2(n14259), .B1(n17939), .B2(n17938), .O(n17941) );
  NR2 U20537 ( .I1(n17942), .I2(n17941), .O(n17943) );
  ND3P U20538 ( .I1(n17945), .I2(n17944), .I3(n17943), .O(n21655) );
  MXL2HS U20539 ( .A(n20863), .B(n21655), .S(n21654), .OB(n20757) );
  INV2 U20540 ( .I(n20757), .O(n20740) );
  AOI22S U20541 ( .A1(n20740), .A2(n19603), .B1(n20527), .B2(n19818), .O(
        n17946) );
  ND3P U20542 ( .I1(n17952), .I2(n17951), .I3(n17950), .O(n22062) );
  ND2S U20543 ( .I1(n22062), .I2(n20809), .O(n17953) );
  BUF2 U20544 ( .I(n17953), .O(n21407) );
  AOI22S U20545 ( .A1(n19603), .A2(n20863), .B1(n20509), .B2(n22923), .O(
        n17955) );
  ND2S U20546 ( .I1(n20509), .I2(n19818), .O(n17954) );
  ND2S U20547 ( .I1(n17955), .I2(n17954), .O(n17956) );
  AN2T U20548 ( .I1(n21808), .I2(n20809), .O(n20535) );
  ND2S U20549 ( .I1(n20535), .I2(n13810), .O(n17963) );
  AOI22S U20550 ( .A1(n13814), .A2(n21601), .B1(n17964), .B2(n17963), .O(
        n17966) );
  ND2S U20551 ( .I1(n22054), .I2(n20809), .O(n17965) );
  OAI22S U20552 ( .A1(n17967), .A2(n17966), .B1(n21804), .B2(n17965), .O(
        n17968) );
  AOI22S U20553 ( .A1(n19326), .A2(img[1010]), .B1(n13837), .B2(img[882]), .O(
        n17973) );
  AOI22S U20554 ( .A1(n15506), .A2(img[754]), .B1(n13858), .B2(img[626]), .O(
        n17972) );
  BUF2 U20555 ( .I(n19642), .O(n19388) );
  AOI22S U20556 ( .A1(n19710), .A2(img[498]), .B1(n19388), .B2(img[370]), .O(
        n17971) );
  AOI22S U20557 ( .A1(n13833), .A2(img[242]), .B1(n18832), .B2(img[114]), .O(
        n17970) );
  AN4S U20558 ( .I1(n17973), .I2(n17972), .I3(n17971), .I4(n17970), .O(n17979)
         );
  AOI22S U20559 ( .A1(n13786), .A2(img[2034]), .B1(n13832), .B2(img[1906]), 
        .O(n17977) );
  AOI22S U20560 ( .A1(n17382), .A2(img[1778]), .B1(n19182), .B2(img[1650]), 
        .O(n17976) );
  AOI22S U20561 ( .A1(n17312), .A2(img[1522]), .B1(n19271), .B2(img[1394]), 
        .O(n17975) );
  AOI22S U20562 ( .A1(n13788), .A2(img[1266]), .B1(n13890), .B2(img[1138]), 
        .O(n17974) );
  AN4S U20563 ( .I1(n17977), .I2(n17976), .I3(n17975), .I4(n17974), .O(n17978)
         );
  ND2P U20564 ( .I1(n17979), .I2(n17978), .O(n19903) );
  AOI22S U20565 ( .A1(n19252), .A2(img[946]), .B1(n13797), .B2(img[818]), .O(
        n17983) );
  AOI22S U20566 ( .A1(n13785), .A2(img[690]), .B1(n13855), .B2(img[562]), .O(
        n17982) );
  BUF1 U20567 ( .I(n19710), .O(n19302) );
  BUF2 U20568 ( .I(n19642), .O(n20103) );
  AOI22S U20569 ( .A1(n19302), .A2(img[434]), .B1(n13836), .B2(img[306]), .O(
        n17981) );
  AOI22S U20570 ( .A1(n13803), .A2(img[178]), .B1(n20193), .B2(img[50]), .O(
        n17980) );
  AN4S U20571 ( .I1(n17983), .I2(n17982), .I3(n17981), .I4(n17980), .O(n17989)
         );
  AOI22S U20572 ( .A1(n19215), .A2(img[1970]), .B1(n13832), .B2(img[1842]), 
        .O(n17987) );
  AOI22S U20573 ( .A1(n13874), .A2(img[1714]), .B1(n19182), .B2(img[1586]), 
        .O(n17986) );
  AOI22S U20574 ( .A1(n13783), .A2(img[1458]), .B1(n15800), .B2(img[1330]), 
        .O(n17985) );
  INV1S U20575 ( .I(n16516), .O(n19127) );
  AOI22S U20576 ( .A1(n18946), .A2(img[1202]), .B1(n13861), .B2(img[1074]), 
        .O(n17984) );
  AN4S U20577 ( .I1(n17987), .I2(n17986), .I3(n17985), .I4(n17984), .O(n17988)
         );
  ND2 U20578 ( .I1(n17989), .I2(n17988), .O(n19885) );
  AOI22S U20579 ( .A1(n19903), .A2(n13839), .B1(n17875), .B2(n19885), .O(
        n18054) );
  AOI22S U20580 ( .A1(n19265), .A2(img[1002]), .B1(n13837), .B2(img[874]), .O(
        n17993) );
  AOI22S U20581 ( .A1(n15506), .A2(img[746]), .B1(n19709), .B2(img[618]), .O(
        n17992) );
  AOI22S U20582 ( .A1(n19266), .A2(img[490]), .B1(n13836), .B2(img[362]), .O(
        n17991) );
  AOI22S U20583 ( .A1(n18797), .A2(img[234]), .B1(n20193), .B2(img[106]), .O(
        n17990) );
  AN4S U20584 ( .I1(n17993), .I2(n17992), .I3(n17991), .I4(n17990), .O(n17999)
         );
  AOI22S U20585 ( .A1(n13786), .A2(img[2026]), .B1(n18201), .B2(img[1898]), 
        .O(n17997) );
  AOI22S U20586 ( .A1(n15630), .A2(img[1770]), .B1(n19182), .B2(img[1642]), 
        .O(n17996) );
  AOI22S U20587 ( .A1(n17359), .A2(img[1514]), .B1(n19271), .B2(img[1386]), 
        .O(n17995) );
  AOI22S U20588 ( .A1(n16515), .A2(img[1258]), .B1(n13890), .B2(img[1130]), 
        .O(n17994) );
  AN4S U20589 ( .I1(n17997), .I2(n17996), .I3(n17995), .I4(n17994), .O(n17998)
         );
  ND2 U20590 ( .I1(n17999), .I2(n17998), .O(n19893) );
  AOI22S U20591 ( .A1(n19252), .A2(img[954]), .B1(n13797), .B2(img[826]), .O(
        n18003) );
  AOI22S U20592 ( .A1(n15506), .A2(img[698]), .B1(n19709), .B2(img[570]), .O(
        n18002) );
  AOI22S U20593 ( .A1(n19253), .A2(img[442]), .B1(n13836), .B2(img[314]), .O(
        n18001) );
  AOI22S U20594 ( .A1(n18773), .A2(img[186]), .B1(n20193), .B2(img[58]), .O(
        n18000) );
  AN4S U20595 ( .I1(n18003), .I2(n18002), .I3(n18001), .I4(n18000), .O(n18009)
         );
  AOI22S U20596 ( .A1(n13786), .A2(img[1978]), .B1(n18201), .B2(img[1850]), 
        .O(n18007) );
  AOI22S U20597 ( .A1(n17382), .A2(img[1722]), .B1(n19182), .B2(img[1594]), 
        .O(n18006) );
  AOI22S U20598 ( .A1(n17312), .A2(img[1466]), .B1(n13792), .B2(img[1338]), 
        .O(n18005) );
  AOI22S U20599 ( .A1(n16037), .A2(img[1210]), .B1(n13861), .B2(img[1082]), 
        .O(n18004) );
  AN4S U20600 ( .I1(n18007), .I2(n18006), .I3(n18005), .I4(n18004), .O(n18008)
         );
  ND2S U20601 ( .I1(n18009), .I2(n18008), .O(n19892) );
  AOI22S U20602 ( .A1(n19893), .A2(n19483), .B1(n20187), .B2(n19892), .O(
        n18053) );
  AOI22S U20603 ( .A1(n19288), .A2(img[962]), .B1(n13837), .B2(img[834]), .O(
        n18013) );
  AOI22S U20604 ( .A1(n20032), .A2(img[706]), .B1(n13855), .B2(img[578]), .O(
        n18012) );
  AOI22S U20605 ( .A1(n19289), .A2(img[450]), .B1(n13836), .B2(img[322]), .O(
        n18011) );
  AOI22S U20606 ( .A1(n13803), .A2(img[194]), .B1(n20193), .B2(img[66]), .O(
        n18010) );
  AN4S U20607 ( .I1(n18013), .I2(n18012), .I3(n18011), .I4(n18010), .O(n18019)
         );
  AOI22S U20608 ( .A1(n19215), .A2(img[1986]), .B1(n18201), .B2(img[1858]), 
        .O(n18017) );
  AOI22S U20609 ( .A1(n19193), .A2(img[1730]), .B1(n19001), .B2(img[1602]), 
        .O(n18016) );
  AOI22S U20610 ( .A1(n17359), .A2(img[1474]), .B1(n19295), .B2(img[1346]), 
        .O(n18015) );
  AOI22S U20611 ( .A1(n13788), .A2(img[1218]), .B1(n13861), .B2(img[1090]), 
        .O(n18014) );
  AOI22S U20612 ( .A1(n19326), .A2(img[938]), .B1(n13898), .B2(img[810]), .O(
        n18023) );
  AOI22S U20613 ( .A1(n13785), .A2(img[682]), .B1(n13855), .B2(img[554]), .O(
        n18022) );
  AOI22S U20614 ( .A1(n19302), .A2(img[426]), .B1(n13836), .B2(img[298]), .O(
        n18021) );
  AOI22S U20615 ( .A1(n13801), .A2(img[170]), .B1(n20193), .B2(img[42]), .O(
        n18020) );
  AN4S U20616 ( .I1(n18023), .I2(n18022), .I3(n18021), .I4(n18020), .O(n18029)
         );
  AOI22S U20617 ( .A1(n19036), .A2(img[1962]), .B1(n18201), .B2(img[1834]), 
        .O(n18027) );
  AOI22S U20618 ( .A1(n17382), .A2(img[1706]), .B1(n18751), .B2(img[1578]), 
        .O(n18026) );
  AOI22S U20619 ( .A1(n16635), .A2(img[1450]), .B1(n20198), .B2(img[1322]), 
        .O(n18025) );
  AOI22S U20620 ( .A1(n16515), .A2(img[1194]), .B1(n13893), .B2(img[1066]), 
        .O(n18024) );
  AN4S U20621 ( .I1(n18027), .I2(n18026), .I3(n18025), .I4(n18024), .O(n18028)
         );
  AOI22S U20622 ( .A1(n19891), .A2(n13843), .B1(n20124), .B2(n19882), .O(
        n18052) );
  AOI22S U20623 ( .A1(n19641), .A2(img[970]), .B1(n13797), .B2(img[842]), .O(
        n18033) );
  AOI22S U20624 ( .A1(n13785), .A2(img[714]), .B1(n13896), .B2(img[586]), .O(
        n18032) );
  AOI22S U20625 ( .A1(n19313), .A2(img[458]), .B1(n13836), .B2(img[330]), .O(
        n18031) );
  AOI22S U20626 ( .A1(n13801), .A2(img[202]), .B1(n20193), .B2(img[74]), .O(
        n18030) );
  AN4S U20627 ( .I1(n18033), .I2(n18032), .I3(n18031), .I4(n18030), .O(n18039)
         );
  AOI22S U20628 ( .A1(n13786), .A2(img[1994]), .B1(n18201), .B2(img[1866]), 
        .O(n18037) );
  AOI22S U20629 ( .A1(n20109), .A2(img[1738]), .B1(n19182), .B2(img[1610]), 
        .O(n18036) );
  AOI22S U20630 ( .A1(n13783), .A2(img[1482]), .B1(n19319), .B2(img[1354]), 
        .O(n18035) );
  AOI22S U20631 ( .A1(n18148), .A2(img[1226]), .B1(n13861), .B2(img[1098]), 
        .O(n18034) );
  AN4S U20632 ( .I1(n18037), .I2(n18036), .I3(n18035), .I4(n18034), .O(n18038)
         );
  ND2 U20633 ( .I1(n18039), .I2(n18038), .O(n19895) );
  AOI22S U20634 ( .A1(n19326), .A2(img[914]), .B1(n13898), .B2(img[786]), .O(
        n18044) );
  AOI22S U20635 ( .A1(n13825), .A2(img[658]), .B1(n13858), .B2(img[530]), .O(
        n18043) );
  BUF1 U20636 ( .I(n19710), .O(n19327) );
  AOI22S U20637 ( .A1(n19327), .A2(img[402]), .B1(n13836), .B2(img[274]), .O(
        n18042) );
  AOI22S U20638 ( .A1(n17335), .A2(img[146]), .B1(n20193), .B2(img[18]), .O(
        n18041) );
  AN4S U20639 ( .I1(n18044), .I2(n18043), .I3(n18042), .I4(n18041), .O(n18050)
         );
  AOI22S U20640 ( .A1(n13786), .A2(img[1938]), .B1(n19416), .B2(img[1810]), 
        .O(n18048) );
  AOI22S U20641 ( .A1(n20109), .A2(img[1682]), .B1(n19182), .B2(img[1554]), 
        .O(n18047) );
  AOI22S U20642 ( .A1(n17336), .A2(img[1426]), .B1(n19319), .B2(img[1298]), 
        .O(n18046) );
  AOI22S U20643 ( .A1(n17810), .A2(img[1170]), .B1(n13893), .B2(img[1042]), 
        .O(n18045) );
  AN4S U20644 ( .I1(n18048), .I2(n18047), .I3(n18046), .I4(n18045), .O(n18049)
         );
  ND2 U20645 ( .I1(n18050), .I2(n18049), .O(n19894) );
  AOI22S U20646 ( .A1(n19895), .A2(n20968), .B1(n13830), .B2(n19894), .O(
        n18051) );
  AN4 U20647 ( .I1(n18054), .I2(n18053), .I3(n18052), .I4(n18051), .O(n18131)
         );
  AOI22S U20648 ( .A1(n19641), .A2(img[978]), .B1(n13837), .B2(img[850]), .O(
        n18058) );
  AOI22S U20649 ( .A1(n15506), .A2(img[722]), .B1(n13855), .B2(img[594]), .O(
        n18057) );
  AOI22S U20650 ( .A1(n19313), .A2(img[466]), .B1(n13836), .B2(img[338]), .O(
        n18056) );
  AOI22S U20651 ( .A1(n17816), .A2(img[210]), .B1(n20193), .B2(img[82]), .O(
        n18055) );
  AN4S U20652 ( .I1(n18058), .I2(n18057), .I3(n18056), .I4(n18055), .O(n18064)
         );
  AOI22S U20653 ( .A1(n19036), .A2(img[2002]), .B1(n17561), .B2(img[1874]), 
        .O(n18062) );
  AOI22S U20654 ( .A1(n17382), .A2(img[1746]), .B1(n13799), .B2(img[1618]), 
        .O(n18061) );
  AOI22S U20655 ( .A1(n13783), .A2(img[1490]), .B1(n19319), .B2(img[1362]), 
        .O(n18060) );
  AOI22S U20656 ( .A1(n13788), .A2(img[1234]), .B1(n16048), .B2(img[1106]), 
        .O(n18059) );
  AOI22S U20657 ( .A1(n19265), .A2(img[906]), .B1(n13898), .B2(img[778]), .O(
        n18068) );
  AOI22S U20658 ( .A1(n13785), .A2(img[650]), .B1(n13855), .B2(img[522]), .O(
        n18067) );
  BUF1 U20659 ( .I(n19710), .O(n20192) );
  AOI22S U20660 ( .A1(n20192), .A2(img[394]), .B1(n13836), .B2(img[266]), .O(
        n18066) );
  AOI22S U20661 ( .A1(n18958), .A2(img[138]), .B1(n20193), .B2(img[10]), .O(
        n18065) );
  AN4S U20662 ( .I1(n18068), .I2(n18067), .I3(n18066), .I4(n18065), .O(n18074)
         );
  AOI22S U20663 ( .A1(n19036), .A2(img[1930]), .B1(n17550), .B2(img[1802]), 
        .O(n18072) );
  AOI22S U20664 ( .A1(n19193), .A2(img[1674]), .B1(n13799), .B2(img[1546]), 
        .O(n18071) );
  AOI22S U20665 ( .A1(n17336), .A2(img[1418]), .B1(n20198), .B2(img[1290]), 
        .O(n18070) );
  AOI22S U20666 ( .A1(n19037), .A2(img[1162]), .B1(n13890), .B2(img[1034]), 
        .O(n18069) );
  AN4S U20667 ( .I1(n18072), .I2(n18071), .I3(n18070), .I4(n18069), .O(n18073)
         );
  ND2 U20668 ( .I1(n18074), .I2(n18073), .O(n19883) );
  AOI22S U20669 ( .A1(n19896), .A2(n20439), .B1(n13847), .B2(n19883), .O(
        n18129) );
  AOI22S U20670 ( .A1(n19326), .A2(img[922]), .B1(n13837), .B2(img[794]), .O(
        n18078) );
  AOI22S U20671 ( .A1(n13825), .A2(img[666]), .B1(n13858), .B2(img[538]), .O(
        n18077) );
  AOI22S U20672 ( .A1(n19327), .A2(img[410]), .B1(n13836), .B2(img[282]), .O(
        n18076) );
  AOI22S U20673 ( .A1(n19290), .A2(img[154]), .B1(n20193), .B2(img[26]), .O(
        n18075) );
  AN4S U20674 ( .I1(n18078), .I2(n18077), .I3(n18076), .I4(n18075), .O(n18084)
         );
  AOI22S U20675 ( .A1(n19215), .A2(img[1946]), .B1(n13794), .B2(img[1818]), 
        .O(n18082) );
  AOI22S U20676 ( .A1(n18837), .A2(img[1690]), .B1(n17827), .B2(img[1562]), 
        .O(n18081) );
  AOI22S U20677 ( .A1(n17347), .A2(img[1434]), .B1(n15800), .B2(img[1306]), 
        .O(n18080) );
  AOI22S U20678 ( .A1(n13788), .A2(img[1178]), .B1(n13877), .B2(img[1050]), 
        .O(n18079) );
  AN4S U20679 ( .I1(n18082), .I2(n18081), .I3(n18080), .I4(n18079), .O(n18083)
         );
  ND2S U20680 ( .I1(n18084), .I2(n18083), .O(n19884) );
  ND2S U20681 ( .I1(n19884), .I2(n17762), .O(n18128) );
  AOI22S U20682 ( .A1(n19376), .A2(img[930]), .B1(n13837), .B2(img[802]), .O(
        n18088) );
  AOI22S U20683 ( .A1(n18681), .A2(img[674]), .B1(n13859), .B2(img[546]), .O(
        n18087) );
  BUF1 U20684 ( .I(n19710), .O(n19377) );
  AOI22S U20685 ( .A1(n19377), .A2(img[418]), .B1(n13836), .B2(img[290]), .O(
        n18086) );
  AOI22S U20686 ( .A1(n18983), .A2(img[162]), .B1(n20193), .B2(img[34]), .O(
        n18085) );
  AN4S U20687 ( .I1(n18088), .I2(n18087), .I3(n18086), .I4(n18085), .O(n18094)
         );
  AOI22S U20688 ( .A1(n13786), .A2(img[1954]), .B1(n17550), .B2(img[1826]), 
        .O(n18092) );
  AOI22S U20689 ( .A1(n19193), .A2(img[1698]), .B1(n17862), .B2(img[1570]), 
        .O(n18091) );
  AOI22S U20690 ( .A1(n17347), .A2(img[1442]), .B1(n13787), .B2(img[1314]), 
        .O(n18090) );
  AOI22S U20691 ( .A1(n16515), .A2(img[1186]), .B1(n13890), .B2(img[1058]), 
        .O(n18089) );
  AN4S U20692 ( .I1(n18092), .I2(n18091), .I3(n18090), .I4(n18089), .O(n18093)
         );
  AOI22S U20693 ( .A1(n19710), .A2(img[506]), .B1(n19388), .B2(img[378]), .O(
        n18098) );
  AOI22S U20694 ( .A1(n13841), .A2(img[250]), .B1(n18832), .B2(img[122]), .O(
        n18097) );
  AOI22S U20695 ( .A1(n19288), .A2(img[1018]), .B1(n13797), .B2(img[890]), .O(
        n18096) );
  AOI22S U20696 ( .A1(n20032), .A2(img[762]), .B1(n15799), .B2(img[634]), .O(
        n18095) );
  AN4S U20697 ( .I1(n18098), .I2(n18097), .I3(n18096), .I4(n18095), .O(n18104)
         );
  AOI22S U20698 ( .A1(n13786), .A2(img[2042]), .B1(n19416), .B2(img[1914]), 
        .O(n18102) );
  AOI22S U20699 ( .A1(n19193), .A2(img[1786]), .B1(n17862), .B2(img[1658]), 
        .O(n18101) );
  AOI22S U20700 ( .A1(n13854), .A2(img[1530]), .B1(n19955), .B2(img[1402]), 
        .O(n18100) );
  AOI22S U20701 ( .A1(n18935), .A2(img[1274]), .B1(n13889), .B2(img[1146]), 
        .O(n18099) );
  AN4S U20702 ( .I1(n18102), .I2(n18101), .I3(n18100), .I4(n18099), .O(n18103)
         );
  AOI22S U20703 ( .A1(n19879), .A2(n13804), .B1(n13846), .B2(n20334), .O(
        n18127) );
  AOI22S U20704 ( .A1(n19342), .A2(img[986]), .B1(n13797), .B2(img[858]), .O(
        n18108) );
  AOI22S U20705 ( .A1(n20102), .A2(img[730]), .B1(n13879), .B2(img[602]), .O(
        n18107) );
  BUF1 U20706 ( .I(n19710), .O(n19344) );
  AOI22S U20707 ( .A1(n19344), .A2(img[474]), .B1(n13836), .B2(img[346]), .O(
        n18106) );
  AOI22S U20708 ( .A1(n14909), .A2(img[218]), .B1(n20193), .B2(img[90]), .O(
        n18105) );
  AN4S U20709 ( .I1(n18108), .I2(n18107), .I3(n18106), .I4(n18105), .O(n18115)
         );
  AOI22S U20710 ( .A1(n19215), .A2(img[2010]), .B1(n18201), .B2(img[1882]), 
        .O(n18113) );
  AOI22S U20711 ( .A1(n19193), .A2(img[1754]), .B1(n17827), .B2(img[1626]), 
        .O(n18112) );
  AOI22S U20712 ( .A1(n13783), .A2(img[1498]), .B1(n19349), .B2(img[1370]), 
        .O(n18111) );
  AOI22S U20713 ( .A1(n18946), .A2(img[1242]), .B1(n15653), .B2(img[1114]), 
        .O(n18110) );
  AN4S U20714 ( .I1(n18113), .I2(n18112), .I3(n18111), .I4(n18110), .O(n18114)
         );
  ND2S U20715 ( .I1(n18115), .I2(n18114), .O(n19881) );
  AOI22S U20716 ( .A1(n19288), .A2(img[994]), .B1(n13837), .B2(img[866]), .O(
        n18119) );
  AOI22S U20717 ( .A1(n13785), .A2(img[738]), .B1(n13896), .B2(img[610]), .O(
        n18118) );
  BUF1 U20718 ( .I(n19710), .O(n19410) );
  AOI22S U20719 ( .A1(n19410), .A2(img[482]), .B1(n13836), .B2(img[354]), .O(
        n18117) );
  AOI22S U20720 ( .A1(n18819), .A2(img[226]), .B1(n20193), .B2(img[98]), .O(
        n18116) );
  AN4S U20721 ( .I1(n18119), .I2(n18118), .I3(n18117), .I4(n18116), .O(n18125)
         );
  AOI22S U20722 ( .A1(n13786), .A2(img[2018]), .B1(n18201), .B2(img[1890]), 
        .O(n18123) );
  AOI22S U20723 ( .A1(n19193), .A2(img[1762]), .B1(n17827), .B2(img[1634]), 
        .O(n18122) );
  AOI22S U20724 ( .A1(n17088), .A2(img[1506]), .B1(n19417), .B2(img[1378]), 
        .O(n18121) );
  AOI22S U20725 ( .A1(n20110), .A2(img[1250]), .B1(n13890), .B2(img[1122]), 
        .O(n18120) );
  ND2S U20726 ( .I1(n18125), .I2(n18124), .O(n19880) );
  AOI22S U20727 ( .A1(n19881), .A2(n13791), .B1(n13835), .B2(n19880), .O(
        n18126) );
  AN4 U20728 ( .I1(n18129), .I2(n18128), .I3(n18127), .I4(n18126), .O(n18130)
         );
  ND2P U20729 ( .I1(n18131), .I2(n18130), .O(n18137) );
  INV1S U20730 ( .I(n18137), .O(n18140) );
  AOI22S U20731 ( .A1(n18137), .A2(n20364), .B1(n20363), .B2(n18137), .O(
        n18139) );
  INV1S U20732 ( .I(n20334), .O(n18135) );
  NR2T U20733 ( .I1(n18134), .I2(n18133), .O(n19600) );
  INV1S U20734 ( .I(n19600), .O(n19430) );
  MOAI1S U20735 ( .A1(n18135), .A2(n19430), .B1(n20334), .B2(n19601), .O(
        n18136) );
  AOI12HS U20736 ( .B1(n18137), .B2(n20373), .A1(n18136), .O(n18138) );
  OAI112HS U20737 ( .C1(n18140), .C2(n19542), .A1(n18139), .B1(n18138), .O(
        n22933) );
  ND2S U20738 ( .I1(n22933), .I2(n20809), .O(n18143) );
  ND2S U20739 ( .I1(n19534), .I2(n18142), .O(n22934) );
  INV1S U20740 ( .I(n29497), .O(n25395) );
  AOI22S U20741 ( .A1(n17835), .A2(img[1011]), .B1(n13797), .B2(img[883]), .O(
        n18147) );
  AOI22S U20742 ( .A1(n20032), .A2(img[755]), .B1(n13858), .B2(img[627]), .O(
        n18146) );
  AOI22S U20743 ( .A1(n19710), .A2(img[499]), .B1(n19388), .B2(img[371]), .O(
        n18145) );
  AOI22S U20744 ( .A1(n13833), .A2(img[243]), .B1(n18832), .B2(img[115]), .O(
        n18144) );
  AN4S U20745 ( .I1(n18147), .I2(n18146), .I3(n18145), .I4(n18144), .O(n18154)
         );
  AOI22S U20746 ( .A1(n18885), .A2(img[2035]), .B1(n18201), .B2(img[1907]), 
        .O(n18152) );
  AOI22S U20747 ( .A1(n19193), .A2(img[1779]), .B1(n13845), .B2(img[1651]), 
        .O(n18151) );
  AOI22S U20748 ( .A1(n18897), .A2(img[1523]), .B1(n20039), .B2(img[1395]), 
        .O(n18150) );
  AOI22S U20749 ( .A1(n16037), .A2(img[1267]), .B1(n13890), .B2(img[1139]), 
        .O(n18149) );
  AN4S U20750 ( .I1(n18152), .I2(n18151), .I3(n18150), .I4(n18149), .O(n18153)
         );
  ND2P U20751 ( .I1(n18154), .I2(n18153), .O(n19701) );
  AOI22S U20752 ( .A1(n13875), .A2(img[947]), .B1(n13837), .B2(img[819]), .O(
        n18159) );
  AOI22S U20753 ( .A1(n18681), .A2(img[691]), .B1(n15799), .B2(img[563]), .O(
        n18158) );
  AOI22S U20754 ( .A1(n19710), .A2(img[435]), .B1(n17611), .B2(img[307]), .O(
        n18157) );
  BUF4 U20755 ( .I(n15080), .O(n19950) );
  AOI22S U20756 ( .A1(n13801), .A2(img[179]), .B1(n19950), .B2(img[51]), .O(
        n18156) );
  AN4S U20757 ( .I1(n18159), .I2(n18158), .I3(n18157), .I4(n18156), .O(n18165)
         );
  AOI22S U20758 ( .A1(n13786), .A2(img[1971]), .B1(n19416), .B2(img[1843]), 
        .O(n18163) );
  AOI22S U20759 ( .A1(n13874), .A2(img[1715]), .B1(n17862), .B2(img[1587]), 
        .O(n18162) );
  INV1S U20760 ( .I(n13789), .O(n18923) );
  AOI22S U20761 ( .A1(n18923), .A2(img[1459]), .B1(n18922), .B2(img[1331]), 
        .O(n18161) );
  AOI22S U20762 ( .A1(n18946), .A2(img[1203]), .B1(n16048), .B2(img[1075]), 
        .O(n18160) );
  ND2 U20763 ( .I1(n18165), .I2(n18164), .O(n19667) );
  AOI22S U20764 ( .A1(n19701), .A2(n13839), .B1(n17875), .B2(n19667), .O(
        n18231) );
  AOI22S U20765 ( .A1(n19326), .A2(img[1003]), .B1(n13837), .B2(img[875]), .O(
        n18169) );
  AOI22S U20766 ( .A1(n18681), .A2(img[747]), .B1(n19709), .B2(img[619]), .O(
        n18168) );
  AOI22S U20767 ( .A1(n19031), .A2(img[491]), .B1(n17611), .B2(img[363]), .O(
        n18167) );
  AOI22S U20768 ( .A1(n18797), .A2(img[235]), .B1(n19950), .B2(img[107]), .O(
        n18166) );
  AOI22S U20769 ( .A1(n19215), .A2(img[2027]), .B1(n13794), .B2(img[1899]), 
        .O(n18173) );
  AOI22S U20770 ( .A1(n13874), .A2(img[1771]), .B1(n13845), .B2(img[1643]), 
        .O(n18172) );
  AOI22S U20771 ( .A1(n18910), .A2(img[1515]), .B1(n13802), .B2(img[1387]), 
        .O(n18171) );
  AOI22S U20772 ( .A1(n16037), .A2(img[1259]), .B1(n16048), .B2(img[1131]), 
        .O(n18170) );
  AN4S U20773 ( .I1(n18173), .I2(n18172), .I3(n18171), .I4(n18170), .O(n18174)
         );
  AOI22S U20774 ( .A1(n19326), .A2(img[955]), .B1(n13837), .B2(img[827]), .O(
        n18179) );
  AOI22S U20775 ( .A1(n13785), .A2(img[699]), .B1(n13855), .B2(img[571]), .O(
        n18178) );
  AOI22S U20776 ( .A1(n18892), .A2(img[443]), .B1(n17611), .B2(img[315]), .O(
        n18177) );
  AOI22S U20777 ( .A1(n13833), .A2(img[187]), .B1(n19950), .B2(img[59]), .O(
        n18176) );
  AN4 U20778 ( .I1(n18179), .I2(n18178), .I3(n18177), .I4(n18176), .O(n18185)
         );
  AOI22S U20779 ( .A1(n13823), .A2(img[1723]), .B1(n13799), .B2(img[1595]), 
        .O(n18182) );
  INV1S U20780 ( .I(n13789), .O(n18897) );
  AOI22S U20781 ( .A1(n18897), .A2(img[1467]), .B1(n18922), .B2(img[1339]), 
        .O(n18181) );
  AOI22S U20782 ( .A1(n20110), .A2(img[1211]), .B1(n13893), .B2(img[1083]), 
        .O(n18180) );
  AOI22S U20783 ( .A1(n19684), .A2(n19483), .B1(n20187), .B2(n19674), .O(
        n18230) );
  AOI22S U20784 ( .A1(n19326), .A2(img[963]), .B1(n13837), .B2(img[835]), .O(
        n18189) );
  AOI22S U20785 ( .A1(n19343), .A2(img[707]), .B1(n13879), .B2(img[579]), .O(
        n18188) );
  BUF1 U20786 ( .I(n19710), .O(n18904) );
  AOI22S U20787 ( .A1(n18904), .A2(img[451]), .B1(n17611), .B2(img[323]), .O(
        n18187) );
  AOI22S U20788 ( .A1(n13841), .A2(img[195]), .B1(n19950), .B2(img[67]), .O(
        n18186) );
  AN4S U20789 ( .I1(n18189), .I2(n18188), .I3(n18187), .I4(n18186), .O(n18195)
         );
  AOI22S U20790 ( .A1(n19036), .A2(img[1987]), .B1(n13832), .B2(img[1859]), 
        .O(n18193) );
  AOI22S U20791 ( .A1(n13874), .A2(img[1731]), .B1(n19182), .B2(img[1603]), 
        .O(n18192) );
  INV1S U20792 ( .I(n13789), .O(n18910) );
  BUF1S U20793 ( .I(n15561), .O(n18909) );
  AOI22S U20794 ( .A1(n18910), .A2(img[1475]), .B1(n18909), .B2(img[1347]), 
        .O(n18191) );
  AOI22S U20795 ( .A1(n19956), .A2(img[1219]), .B1(n15653), .B2(img[1091]), 
        .O(n18190) );
  AN4S U20796 ( .I1(n18193), .I2(n18192), .I3(n18191), .I4(n18190), .O(n18194)
         );
  ND2 U20797 ( .I1(n18195), .I2(n18194), .O(n19673) );
  AOI22S U20798 ( .A1(n13875), .A2(img[939]), .B1(n13837), .B2(img[811]), .O(
        n18200) );
  AOI22S U20799 ( .A1(n13785), .A2(img[683]), .B1(n15691), .B2(img[555]), .O(
        n18199) );
  AOI22S U20800 ( .A1(n19710), .A2(img[427]), .B1(n17611), .B2(img[299]), .O(
        n18198) );
  AOI22S U20801 ( .A1(n14909), .A2(img[171]), .B1(n19950), .B2(img[43]), .O(
        n18197) );
  AN4S U20802 ( .I1(n18200), .I2(n18199), .I3(n18198), .I4(n18197), .O(n18207)
         );
  AOI22S U20803 ( .A1(n19023), .A2(img[1963]), .B1(n18201), .B2(img[1835]), 
        .O(n18205) );
  AOI22S U20804 ( .A1(n13823), .A2(img[1707]), .B1(n19182), .B2(img[1579]), 
        .O(n18204) );
  AOI22S U20805 ( .A1(n18897), .A2(img[1451]), .B1(n18922), .B2(img[1323]), 
        .O(n18203) );
  AOI22S U20806 ( .A1(n14189), .A2(img[1195]), .B1(n15653), .B2(img[1067]), 
        .O(n18202) );
  ND2P U20807 ( .I1(n18207), .I2(n18206), .O(n19685) );
  AOI22S U20808 ( .A1(n19673), .A2(n13843), .B1(n20124), .B2(n19685), .O(
        n18229) );
  AOI22S U20809 ( .A1(n19326), .A2(img[971]), .B1(n13837), .B2(img[843]), .O(
        n18211) );
  AOI22S U20810 ( .A1(n15506), .A2(img[715]), .B1(n13858), .B2(img[587]), .O(
        n18210) );
  AOI22S U20811 ( .A1(n18904), .A2(img[459]), .B1(n17611), .B2(img[331]), .O(
        n18209) );
  AOI22S U20812 ( .A1(n19290), .A2(img[203]), .B1(n19950), .B2(img[75]), .O(
        n18208) );
  AN4S U20813 ( .I1(n18211), .I2(n18210), .I3(n18209), .I4(n18208), .O(n18217)
         );
  AOI22S U20814 ( .A1(n19023), .A2(img[1995]), .B1(n18201), .B2(img[1867]), 
        .O(n18215) );
  AOI22S U20815 ( .A1(n18837), .A2(img[1739]), .B1(n19001), .B2(img[1611]), 
        .O(n18214) );
  AOI22S U20816 ( .A1(n18910), .A2(img[1483]), .B1(n18909), .B2(img[1355]), 
        .O(n18213) );
  AOI22S U20817 ( .A1(n19037), .A2(img[1227]), .B1(n13893), .B2(img[1099]), 
        .O(n18212) );
  AOI22S U20818 ( .A1(n13875), .A2(img[915]), .B1(n13797), .B2(img[787]), .O(
        n18221) );
  AOI22S U20819 ( .A1(n15506), .A2(img[659]), .B1(n13859), .B2(img[531]), .O(
        n18220) );
  AOI22S U20820 ( .A1(n19710), .A2(img[403]), .B1(n17611), .B2(img[275]), .O(
        n18219) );
  AOI22S U20821 ( .A1(n13841), .A2(img[147]), .B1(n19950), .B2(img[19]), .O(
        n18218) );
  AN4S U20822 ( .I1(n18221), .I2(n18220), .I3(n18219), .I4(n18218), .O(n18227)
         );
  AOI22S U20823 ( .A1(n19215), .A2(img[1939]), .B1(n19416), .B2(img[1811]), 
        .O(n18225) );
  BUF1 U20824 ( .I(n13845), .O(n19001) );
  AOI22S U20825 ( .A1(n19193), .A2(img[1683]), .B1(n19001), .B2(img[1555]), 
        .O(n18224) );
  INV1S U20826 ( .I(n13789), .O(n19856) );
  AOI22S U20827 ( .A1(n19856), .A2(img[1427]), .B1(n18974), .B2(img[1299]), 
        .O(n18223) );
  AOI22S U20828 ( .A1(n18911), .A2(img[1171]), .B1(n13892), .B2(img[1043]), 
        .O(n18222) );
  AN4S U20829 ( .I1(n18225), .I2(n18224), .I3(n18223), .I4(n18222), .O(n18226)
         );
  ND2 U20830 ( .I1(n18227), .I2(n18226), .O(n19675) );
  AOI22S U20831 ( .A1(n19677), .A2(n20560), .B1(n13830), .B2(n19675), .O(
        n18228) );
  AN4S U20832 ( .I1(n18231), .I2(n18230), .I3(n18229), .I4(n18228), .O(n18310)
         );
  AOI22S U20833 ( .A1(n19326), .A2(img[979]), .B1(n13797), .B2(img[851]), .O(
        n18235) );
  AOI22S U20834 ( .A1(n13785), .A2(img[723]), .B1(n13859), .B2(img[595]), .O(
        n18234) );
  BUF1 U20835 ( .I(n19710), .O(n18957) );
  AOI22S U20836 ( .A1(n18957), .A2(img[467]), .B1(n17611), .B2(img[339]), .O(
        n18233) );
  AOI22S U20837 ( .A1(n17335), .A2(img[211]), .B1(n19950), .B2(img[83]), .O(
        n18232) );
  AN4S U20838 ( .I1(n18235), .I2(n18234), .I3(n18233), .I4(n18232), .O(n18241)
         );
  AOI22S U20839 ( .A1(n13870), .A2(img[2003]), .B1(n18201), .B2(img[1875]), 
        .O(n18239) );
  AOI22S U20840 ( .A1(n13874), .A2(img[1747]), .B1(n13845), .B2(img[1619]), 
        .O(n18238) );
  INV1S U20841 ( .I(n13789), .O(n18963) );
  AOI22S U20842 ( .A1(n18963), .A2(img[1491]), .B1(n13787), .B2(img[1363]), 
        .O(n18237) );
  AOI22S U20843 ( .A1(n18988), .A2(img[1235]), .B1(n13889), .B2(img[1107]), 
        .O(n18236) );
  AN4S U20844 ( .I1(n18239), .I2(n18238), .I3(n18237), .I4(n18236), .O(n18240)
         );
  ND2 U20845 ( .I1(n18241), .I2(n18240), .O(n19676) );
  AOI22S U20846 ( .A1(n19326), .A2(img[907]), .B1(n13837), .B2(img[779]), .O(
        n18245) );
  AOI22S U20847 ( .A1(n18681), .A2(img[651]), .B1(n13858), .B2(img[523]), .O(
        n18244) );
  AOI22S U20848 ( .A1(n19710), .A2(img[395]), .B1(n17611), .B2(img[267]), .O(
        n18243) );
  AOI22S U20849 ( .A1(n18996), .A2(img[139]), .B1(n19950), .B2(img[11]), .O(
        n18242) );
  AOI22S U20850 ( .A1(n13786), .A2(img[1931]), .B1(n17550), .B2(img[1803]), 
        .O(n18249) );
  AOI22S U20851 ( .A1(n19193), .A2(img[1675]), .B1(n17862), .B2(img[1547]), 
        .O(n18248) );
  AOI22S U20852 ( .A1(n18923), .A2(img[1419]), .B1(n18974), .B2(img[1291]), 
        .O(n18247) );
  AOI22S U20853 ( .A1(n19649), .A2(img[1163]), .B1(n13861), .B2(img[1035]), 
        .O(n18246) );
  AN4S U20854 ( .I1(n18249), .I2(n18248), .I3(n18247), .I4(n18246), .O(n18250)
         );
  ND2 U20855 ( .I1(n18251), .I2(n18250), .O(n19665) );
  AOI22S U20856 ( .A1(n19676), .A2(n20263), .B1(n13847), .B2(n19665), .O(
        n18308) );
  AOI22S U20857 ( .A1(n13875), .A2(img[923]), .B1(n13837), .B2(img[795]), .O(
        n18255) );
  AOI22S U20858 ( .A1(n13785), .A2(img[667]), .B1(n13855), .B2(img[539]), .O(
        n18254) );
  BUF1 U20859 ( .I(n19710), .O(n18982) );
  AOI22S U20860 ( .A1(n18982), .A2(img[411]), .B1(n17611), .B2(img[283]), .O(
        n18253) );
  AOI22S U20861 ( .A1(n13803), .A2(img[155]), .B1(n19950), .B2(img[27]), .O(
        n18252) );
  AN4S U20862 ( .I1(n18255), .I2(n18254), .I3(n18253), .I4(n18252), .O(n18261)
         );
  AOI22S U20863 ( .A1(n19023), .A2(img[1947]), .B1(n13794), .B2(img[1819]), 
        .O(n18259) );
  AOI22S U20864 ( .A1(n15630), .A2(img[1691]), .B1(n19182), .B2(img[1563]), 
        .O(n18258) );
  AOI22S U20865 ( .A1(n13824), .A2(img[1435]), .B1(n17865), .B2(img[1307]), 
        .O(n18257) );
  AOI22S U20866 ( .A1(n19956), .A2(img[1179]), .B1(n13890), .B2(img[1051]), 
        .O(n18256) );
  AN4S U20867 ( .I1(n18259), .I2(n18258), .I3(n18257), .I4(n18256), .O(n18260)
         );
  ND2 U20868 ( .I1(n18261), .I2(n18260), .O(n19666) );
  ND2S U20869 ( .I1(n19666), .I2(n17762), .O(n18307) );
  AOI22S U20870 ( .A1(n13875), .A2(img[931]), .B1(n13797), .B2(img[803]), .O(
        n18266) );
  AOI22S U20871 ( .A1(n18681), .A2(img[675]), .B1(n18262), .B2(img[547]), .O(
        n18265) );
  BUF1 U20872 ( .I(n19710), .O(n18995) );
  AOI22S U20873 ( .A1(n18995), .A2(img[419]), .B1(n17611), .B2(img[291]), .O(
        n18264) );
  AOI22S U20874 ( .A1(n13841), .A2(img[163]), .B1(n19950), .B2(img[35]), .O(
        n18263) );
  AN4S U20875 ( .I1(n18266), .I2(n18265), .I3(n18264), .I4(n18263), .O(n18272)
         );
  AOI22S U20876 ( .A1(n19036), .A2(img[1955]), .B1(n19715), .B2(img[1827]), 
        .O(n18270) );
  AOI22S U20877 ( .A1(n19193), .A2(img[1699]), .B1(n19001), .B2(img[1571]), 
        .O(n18269) );
  AOI22S U20878 ( .A1(n19856), .A2(img[1443]), .B1(n13792), .B2(img[1315]), 
        .O(n18268) );
  AOI22S U20879 ( .A1(n18911), .A2(img[1187]), .B1(n16048), .B2(img[1059]), 
        .O(n18267) );
  AN4S U20880 ( .I1(n18270), .I2(n18269), .I3(n18268), .I4(n18267), .O(n18271)
         );
  ND2 U20881 ( .I1(n18272), .I2(n18271), .O(n19662) );
  AOI22S U20882 ( .A1(n19710), .A2(img[507]), .B1(n19388), .B2(img[379]), .O(
        n18276) );
  AOI22S U20883 ( .A1(n13803), .A2(img[251]), .B1(n18832), .B2(img[123]), .O(
        n18275) );
  AOI22S U20884 ( .A1(n19288), .A2(img[1019]), .B1(n13837), .B2(img[891]), .O(
        n18274) );
  AOI22S U20885 ( .A1(n20032), .A2(img[763]), .B1(n19709), .B2(img[635]), .O(
        n18273) );
  AN4S U20886 ( .I1(n18276), .I2(n18275), .I3(n18274), .I4(n18273), .O(n18282)
         );
  AOI22S U20887 ( .A1(n19215), .A2(img[2043]), .B1(n19416), .B2(img[1915]), 
        .O(n18280) );
  AOI22S U20888 ( .A1(n19193), .A2(img[1787]), .B1(n13798), .B2(img[1659]), 
        .O(n18279) );
  AOI22S U20889 ( .A1(n13854), .A2(img[1531]), .B1(n18922), .B2(img[1403]), 
        .O(n18278) );
  AOI22S U20890 ( .A1(n14822), .A2(img[1275]), .B1(n15653), .B2(img[1147]), 
        .O(n18277) );
  AN4S U20891 ( .I1(n18280), .I2(n18279), .I3(n18278), .I4(n18277), .O(n18281)
         );
  ND2P U20892 ( .I1(n18282), .I2(n18281), .O(n20315) );
  AOI22S U20893 ( .A1(n19662), .A2(n13804), .B1(n13846), .B2(n20315), .O(
        n18306) );
  AOI22S U20894 ( .A1(n19326), .A2(img[987]), .B1(n13797), .B2(img[859]), .O(
        n18286) );
  AOI22S U20895 ( .A1(n19343), .A2(img[731]), .B1(n13858), .B2(img[603]), .O(
        n18285) );
  BUF1 U20896 ( .I(n19710), .O(n19018) );
  AOI22S U20897 ( .A1(n19018), .A2(img[475]), .B1(n17611), .B2(img[347]), .O(
        n18284) );
  AOI22S U20898 ( .A1(n13803), .A2(img[219]), .B1(n19950), .B2(img[91]), .O(
        n18283) );
  AN4S U20899 ( .I1(n18286), .I2(n18285), .I3(n18284), .I4(n18283), .O(n18292)
         );
  AOI22S U20900 ( .A1(n19023), .A2(img[2011]), .B1(n13794), .B2(img[1883]), 
        .O(n18290) );
  AOI22S U20901 ( .A1(n13874), .A2(img[1755]), .B1(n17862), .B2(img[1627]), 
        .O(n18289) );
  AOI22S U20902 ( .A1(n13824), .A2(img[1499]), .B1(n19349), .B2(img[1371]), 
        .O(n18288) );
  AOI22S U20903 ( .A1(n19649), .A2(img[1243]), .B1(n13889), .B2(img[1115]), 
        .O(n18287) );
  ND2 U20904 ( .I1(n18292), .I2(n18291), .O(n19664) );
  AOI22S U20905 ( .A1(n19326), .A2(img[995]), .B1(n13797), .B2(img[867]), .O(
        n18296) );
  AOI22S U20906 ( .A1(n15657), .A2(img[739]), .B1(n13855), .B2(img[611]), .O(
        n18295) );
  AOI22S U20907 ( .A1(n19031), .A2(img[483]), .B1(n17611), .B2(img[355]), .O(
        n18294) );
  AOI22S U20908 ( .A1(n17778), .A2(img[227]), .B1(n19950), .B2(img[99]), .O(
        n18293) );
  AN4S U20909 ( .I1(n18296), .I2(n18295), .I3(n18294), .I4(n18293), .O(n18304)
         );
  AOI22S U20910 ( .A1(n19036), .A2(img[2019]), .B1(n13832), .B2(img[1891]), 
        .O(n18302) );
  AOI22S U20911 ( .A1(n13874), .A2(img[1763]), .B1(n17827), .B2(img[1635]), 
        .O(n18301) );
  AOI22S U20912 ( .A1(n18298), .A2(img[1507]), .B1(n13802), .B2(img[1379]), 
        .O(n18300) );
  AOI22S U20913 ( .A1(n13788), .A2(img[1251]), .B1(n13877), .B2(img[1123]), 
        .O(n18299) );
  AN4S U20914 ( .I1(n18302), .I2(n18301), .I3(n18300), .I4(n18299), .O(n18303)
         );
  AOI22S U20915 ( .A1(n19664), .A2(n13791), .B1(n13835), .B2(n19663), .O(
        n18305) );
  AN4S U20916 ( .I1(n18308), .I2(n18307), .I3(n18306), .I4(n18305), .O(n18309)
         );
  INV1S U20917 ( .I(n18315), .O(n18318) );
  INV1S U20918 ( .I(n20363), .O(n19235) );
  AOI22S U20919 ( .A1(n18315), .A2(n20371), .B1(n20364), .B2(n18315), .O(
        n18317) );
  ND2S U20920 ( .I1(n20315), .I2(n19600), .O(n18313) );
  ND2S U20921 ( .I1(n19601), .I2(n20315), .O(n18312) );
  ND2S U20922 ( .I1(n19514), .I2(n18142), .O(n18311) );
  ND3S U20923 ( .I1(n18313), .I2(n18312), .I3(n18311), .O(n18314) );
  AOI12HS U20924 ( .B1(n18315), .B2(n20373), .A1(n18314), .O(n18316) );
  ND2P U20925 ( .I1(n22931), .I2(n20809), .O(n18319) );
  INV1S U20926 ( .I(n29455), .O(n27266) );
  OAI22S U20927 ( .A1(n25395), .A2(n20644), .B1(n20503), .B2(n27266), .O(
        n18670) );
  AOI22S U20928 ( .A1(n17835), .A2(img[1008]), .B1(n13837), .B2(img[880]), .O(
        n18323) );
  AOI22S U20929 ( .A1(n15506), .A2(img[752]), .B1(n19709), .B2(img[624]), .O(
        n18322) );
  AOI22S U20930 ( .A1(n19710), .A2(img[496]), .B1(n19388), .B2(img[368]), .O(
        n18321) );
  AOI22S U20931 ( .A1(n14909), .A2(img[240]), .B1(n18832), .B2(img[112]), .O(
        n18320) );
  AN4S U20932 ( .I1(n18323), .I2(n18322), .I3(n18321), .I4(n18320), .O(n18329)
         );
  AOI22S U20933 ( .A1(n13786), .A2(img[2032]), .B1(n18201), .B2(img[1904]), 
        .O(n18327) );
  AOI22S U20934 ( .A1(n19193), .A2(img[1776]), .B1(n13799), .B2(img[1648]), 
        .O(n18326) );
  AOI22S U20935 ( .A1(n18789), .A2(img[1520]), .B1(n19271), .B2(img[1392]), 
        .O(n18325) );
  AOI22S U20936 ( .A1(n13788), .A2(img[1264]), .B1(n13889), .B2(img[1136]), 
        .O(n18324) );
  AOI22S U20937 ( .A1(n19342), .A2(img[944]), .B1(n13797), .B2(img[816]), .O(
        n18333) );
  AOI22S U20938 ( .A1(n18681), .A2(img[688]), .B1(n13855), .B2(img[560]), .O(
        n18332) );
  AOI22S U20939 ( .A1(n19302), .A2(img[432]), .B1(n13836), .B2(img[304]), .O(
        n18331) );
  AOI22S U20940 ( .A1(n18819), .A2(img[176]), .B1(n20193), .B2(img[48]), .O(
        n18330) );
  AN4S U20941 ( .I1(n18333), .I2(n18332), .I3(n18331), .I4(n18330), .O(n18339)
         );
  AOI22S U20942 ( .A1(n19036), .A2(img[1968]), .B1(n18201), .B2(img[1840]), 
        .O(n18337) );
  AOI22S U20943 ( .A1(n15630), .A2(img[1712]), .B1(n19182), .B2(img[1584]), 
        .O(n18336) );
  AOI22S U20944 ( .A1(n13853), .A2(img[1456]), .B1(n17840), .B2(img[1328]), 
        .O(n18335) );
  AOI22S U20945 ( .A1(n18946), .A2(img[1200]), .B1(n13861), .B2(img[1072]), 
        .O(n18334) );
  AN4S U20946 ( .I1(n18337), .I2(n18336), .I3(n18335), .I4(n18334), .O(n18338)
         );
  ND2 U20947 ( .I1(n18339), .I2(n18338), .O(n19807) );
  AOI22S U20948 ( .A1(n19837), .A2(n13839), .B1(n17875), .B2(n19807), .O(
        n18361) );
  AOI22S U20949 ( .A1(n19342), .A2(img[1000]), .B1(n13837), .B2(img[872]), .O(
        n18343) );
  AOI22S U20950 ( .A1(n20102), .A2(img[744]), .B1(n19709), .B2(img[616]), .O(
        n18342) );
  AOI22S U20951 ( .A1(n19410), .A2(img[488]), .B1(n13836), .B2(img[360]), .O(
        n18341) );
  AOI22S U20952 ( .A1(n13833), .A2(img[232]), .B1(n20193), .B2(img[104]), .O(
        n18340) );
  AN4S U20953 ( .I1(n18343), .I2(n18342), .I3(n18341), .I4(n18340), .O(n18349)
         );
  AOI22S U20954 ( .A1(n19215), .A2(img[2024]), .B1(n18201), .B2(img[1896]), 
        .O(n18347) );
  AOI22S U20955 ( .A1(n18837), .A2(img[1768]), .B1(n19182), .B2(img[1640]), 
        .O(n18346) );
  AOI22S U20956 ( .A1(n17323), .A2(img[1512]), .B1(n19417), .B2(img[1384]), 
        .O(n18345) );
  AOI22S U20957 ( .A1(n19649), .A2(img[1256]), .B1(n16048), .B2(img[1128]), 
        .O(n18344) );
  AN4S U20958 ( .I1(n18347), .I2(n18346), .I3(n18345), .I4(n18344), .O(n18348)
         );
  AOI22S U20959 ( .A1(n19252), .A2(img[952]), .B1(n13797), .B2(img[824]), .O(
        n18353) );
  AOI22S U20960 ( .A1(n13785), .A2(img[696]), .B1(n13896), .B2(img[568]), .O(
        n18352) );
  AOI22S U20961 ( .A1(n19253), .A2(img[440]), .B1(n13836), .B2(img[312]), .O(
        n18351) );
  AOI22S U20962 ( .A1(n14909), .A2(img[184]), .B1(n20193), .B2(img[56]), .O(
        n18350) );
  AN4S U20963 ( .I1(n18353), .I2(n18352), .I3(n18351), .I4(n18350), .O(n18359)
         );
  AOI22S U20964 ( .A1(n13786), .A2(img[1976]), .B1(n18201), .B2(img[1848]), 
        .O(n18357) );
  AOI22S U20965 ( .A1(n19193), .A2(img[1720]), .B1(n19182), .B2(img[1592]), 
        .O(n18356) );
  AOI22S U20966 ( .A1(n13783), .A2(img[1464]), .B1(n13792), .B2(img[1336]), 
        .O(n18355) );
  AOI22S U20967 ( .A1(n18935), .A2(img[1208]), .B1(n15653), .B2(img[1080]), 
        .O(n18354) );
  AN4S U20968 ( .I1(n18357), .I2(n18356), .I3(n18355), .I4(n18354), .O(n18358)
         );
  AOI22S U20969 ( .A1(n19835), .A2(n19483), .B1(n20187), .B2(n19839), .O(
        n18360) );
  ND2S U20970 ( .I1(n18361), .I2(n18360), .O(n18405) );
  AOI22S U20971 ( .A1(n19288), .A2(img[960]), .B1(n13837), .B2(img[832]), .O(
        n18365) );
  AOI22S U20972 ( .A1(n15506), .A2(img[704]), .B1(n13855), .B2(img[576]), .O(
        n18364) );
  AOI22S U20973 ( .A1(n19289), .A2(img[448]), .B1(n13836), .B2(img[320]), .O(
        n18363) );
  AOI22S U20974 ( .A1(n18983), .A2(img[192]), .B1(n20193), .B2(img[64]), .O(
        n18362) );
  AOI22S U20975 ( .A1(n20109), .A2(img[1728]), .B1(n19182), .B2(img[1600]), 
        .O(n18368) );
  AOI22S U20976 ( .A1(n18975), .A2(img[1472]), .B1(n19295), .B2(img[1344]), 
        .O(n18367) );
  AOI22S U20977 ( .A1(n19649), .A2(img[1216]), .B1(n13890), .B2(img[1088]), 
        .O(n18366) );
  AOI22S U20978 ( .A1(n19265), .A2(img[936]), .B1(n13898), .B2(img[808]), .O(
        n18375) );
  AOI22S U20979 ( .A1(n13825), .A2(img[680]), .B1(n13896), .B2(img[552]), .O(
        n18374) );
  AOI22S U20980 ( .A1(n19302), .A2(img[424]), .B1(n13836), .B2(img[296]), .O(
        n18373) );
  AOI22S U20981 ( .A1(n17793), .A2(img[168]), .B1(n20193), .B2(img[40]), .O(
        n18372) );
  AN4S U20982 ( .I1(n18375), .I2(n18374), .I3(n18373), .I4(n18372), .O(n18381)
         );
  AOI22S U20983 ( .A1(n19036), .A2(img[1960]), .B1(n13832), .B2(img[1832]), 
        .O(n18379) );
  AOI22S U20984 ( .A1(n20109), .A2(img[1704]), .B1(n19182), .B2(img[1576]), 
        .O(n18378) );
  AOI22S U20985 ( .A1(n19856), .A2(img[1448]), .B1(n17276), .B2(img[1320]), 
        .O(n18377) );
  AOI22S U20986 ( .A1(n13788), .A2(img[1192]), .B1(n16048), .B2(img[1064]), 
        .O(n18376) );
  AN4S U20987 ( .I1(n18379), .I2(n18378), .I3(n18377), .I4(n18376), .O(n18380)
         );
  AOI22S U20988 ( .A1(n19833), .A2(n13843), .B1(n20124), .B2(n19827), .O(
        n18403) );
  AOI22S U20989 ( .A1(n19288), .A2(img[968]), .B1(n13898), .B2(img[840]), .O(
        n18385) );
  AOI22S U20990 ( .A1(n15506), .A2(img[712]), .B1(n13858), .B2(img[584]), .O(
        n18384) );
  AOI22S U20991 ( .A1(n19289), .A2(img[456]), .B1(n13836), .B2(img[328]), .O(
        n18383) );
  AOI22S U20992 ( .A1(n17778), .A2(img[200]), .B1(n20193), .B2(img[72]), .O(
        n18382) );
  AN4S U20993 ( .I1(n18385), .I2(n18384), .I3(n18383), .I4(n18382), .O(n18391)
         );
  AOI22S U20994 ( .A1(n13786), .A2(img[1992]), .B1(n18201), .B2(img[1864]), 
        .O(n18389) );
  AOI22S U20995 ( .A1(n19193), .A2(img[1736]), .B1(n19182), .B2(img[1608]), 
        .O(n18388) );
  AOI22S U20996 ( .A1(n17323), .A2(img[1480]), .B1(n19295), .B2(img[1352]), 
        .O(n18387) );
  AOI22S U20997 ( .A1(n14505), .A2(img[1224]), .B1(n13877), .B2(img[1096]), 
        .O(n18386) );
  AN4S U20998 ( .I1(n18389), .I2(n18388), .I3(n18387), .I4(n18386), .O(n18390)
         );
  AOI22S U20999 ( .A1(n18702), .A2(img[912]), .B1(n13797), .B2(img[784]), .O(
        n18395) );
  AOI22S U21000 ( .A1(n18681), .A2(img[656]), .B1(n13858), .B2(img[528]), .O(
        n18394) );
  AOI22S U21001 ( .A1(n20192), .A2(img[400]), .B1(n13836), .B2(img[272]), .O(
        n18393) );
  AOI22S U21002 ( .A1(n13803), .A2(img[144]), .B1(n20193), .B2(img[16]), .O(
        n18392) );
  AN4S U21003 ( .I1(n18395), .I2(n18394), .I3(n18393), .I4(n18392), .O(n18401)
         );
  AOI22S U21004 ( .A1(n19215), .A2(img[1936]), .B1(n19416), .B2(img[1808]), 
        .O(n18399) );
  AOI22S U21005 ( .A1(n15630), .A2(img[1680]), .B1(n17862), .B2(img[1552]), 
        .O(n18398) );
  AOI22S U21006 ( .A1(n13783), .A2(img[1424]), .B1(n20198), .B2(img[1296]), 
        .O(n18397) );
  AOI22S U21007 ( .A1(n18988), .A2(img[1168]), .B1(n13890), .B2(img[1040]), 
        .O(n18396) );
  AN4S U21008 ( .I1(n18399), .I2(n18398), .I3(n18397), .I4(n18396), .O(n18400)
         );
  ND2 U21009 ( .I1(n18401), .I2(n18400), .O(n19840) );
  AOI22S U21010 ( .A1(n19825), .A2(n20560), .B1(n13830), .B2(n19840), .O(
        n18402) );
  ND2 U21011 ( .I1(n18403), .I2(n18402), .O(n18404) );
  NR2 U21012 ( .I1(n18405), .I2(n18404), .O(n18483) );
  AOI22S U21013 ( .A1(n19641), .A2(img[976]), .B1(n13797), .B2(img[848]), .O(
        n18409) );
  AOI22S U21014 ( .A1(n13785), .A2(img[720]), .B1(n19709), .B2(img[592]), .O(
        n18408) );
  AOI22S U21015 ( .A1(n19313), .A2(img[464]), .B1(n13836), .B2(img[336]), .O(
        n18407) );
  AOI22S U21016 ( .A1(n17886), .A2(img[208]), .B1(n20193), .B2(img[80]), .O(
        n18406) );
  AN4S U21017 ( .I1(n18409), .I2(n18408), .I3(n18407), .I4(n18406), .O(n18415)
         );
  AOI22S U21018 ( .A1(n13786), .A2(img[2000]), .B1(n18201), .B2(img[1872]), 
        .O(n18413) );
  AOI22S U21019 ( .A1(n13874), .A2(img[1744]), .B1(n16353), .B2(img[1616]), 
        .O(n18412) );
  AOI22S U21020 ( .A1(n13783), .A2(img[1488]), .B1(n19319), .B2(img[1360]), 
        .O(n18411) );
  AOI22S U21021 ( .A1(n14189), .A2(img[1232]), .B1(n13861), .B2(img[1104]), 
        .O(n18410) );
  AOI22S U21022 ( .A1(n13784), .A2(img[904]), .B1(n13837), .B2(img[776]), .O(
        n18419) );
  AOI22S U21023 ( .A1(n15506), .A2(img[648]), .B1(n13858), .B2(img[520]), .O(
        n18418) );
  AOI22S U21024 ( .A1(n20192), .A2(img[392]), .B1(n13836), .B2(img[264]), .O(
        n18417) );
  AOI22S U21025 ( .A1(n13801), .A2(img[136]), .B1(n20193), .B2(img[8]), .O(
        n18416) );
  AN4S U21026 ( .I1(n18419), .I2(n18418), .I3(n18417), .I4(n18416), .O(n18425)
         );
  AOI22S U21027 ( .A1(n13870), .A2(img[1928]), .B1(n13794), .B2(img[1800]), 
        .O(n18423) );
  AOI22S U21028 ( .A1(n13823), .A2(img[1672]), .B1(n19182), .B2(img[1544]), 
        .O(n18422) );
  AOI22S U21029 ( .A1(n18778), .A2(img[1416]), .B1(n20198), .B2(img[1288]), 
        .O(n18421) );
  AOI22S U21030 ( .A1(n14505), .A2(img[1160]), .B1(n13889), .B2(img[1032]), 
        .O(n18420) );
  AN4S U21031 ( .I1(n18423), .I2(n18422), .I3(n18421), .I4(n18420), .O(n18424)
         );
  AOI22S U21032 ( .A1(n19838), .A2(n20263), .B1(n13847), .B2(n19834), .O(
        n18437) );
  AOI22S U21033 ( .A1(n19326), .A2(img[920]), .B1(n13797), .B2(img[792]), .O(
        n18429) );
  AOI22S U21034 ( .A1(n13825), .A2(img[664]), .B1(n13858), .B2(img[536]), .O(
        n18428) );
  AOI22S U21035 ( .A1(n19327), .A2(img[408]), .B1(n13836), .B2(img[280]), .O(
        n18427) );
  AOI22S U21036 ( .A1(n13803), .A2(img[152]), .B1(n20193), .B2(img[24]), .O(
        n18426) );
  AN4S U21037 ( .I1(n18429), .I2(n18428), .I3(n18427), .I4(n18426), .O(n18435)
         );
  AOI22S U21038 ( .A1(n13786), .A2(img[1944]), .B1(n13794), .B2(img[1816]), 
        .O(n18433) );
  AOI22S U21039 ( .A1(n15630), .A2(img[1688]), .B1(n17862), .B2(img[1560]), 
        .O(n18432) );
  AOI22S U21040 ( .A1(n13853), .A2(img[1432]), .B1(n20198), .B2(img[1304]), 
        .O(n18431) );
  AOI22S U21041 ( .A1(n17810), .A2(img[1176]), .B1(n15653), .B2(img[1048]), 
        .O(n18430) );
  ND2 U21042 ( .I1(n18435), .I2(n18434), .O(n19826) );
  ND2S U21043 ( .I1(n19826), .I2(n17762), .O(n18436) );
  ND2S U21044 ( .I1(n18437), .I2(n18436), .O(n18481) );
  AOI22S U21045 ( .A1(n19376), .A2(img[928]), .B1(n13898), .B2(img[800]), .O(
        n18441) );
  AOI22S U21046 ( .A1(n13825), .A2(img[672]), .B1(n13858), .B2(img[544]), .O(
        n18440) );
  AOI22S U21047 ( .A1(n19377), .A2(img[416]), .B1(n13836), .B2(img[288]), .O(
        n18439) );
  AOI22S U21048 ( .A1(n17864), .A2(img[160]), .B1(n20193), .B2(img[32]), .O(
        n18438) );
  AN4S U21049 ( .I1(n18441), .I2(n18440), .I3(n18439), .I4(n18438), .O(n18447)
         );
  AOI22S U21050 ( .A1(n13786), .A2(img[1952]), .B1(n18201), .B2(img[1824]), 
        .O(n18445) );
  AOI22S U21051 ( .A1(n17382), .A2(img[1696]), .B1(n19182), .B2(img[1568]), 
        .O(n18444) );
  AOI22S U21052 ( .A1(n13853), .A2(img[1440]), .B1(n18623), .B2(img[1312]), 
        .O(n18443) );
  AOI22S U21053 ( .A1(n18148), .A2(img[1184]), .B1(n13890), .B2(img[1056]), 
        .O(n18442) );
  AOI22S U21054 ( .A1(n19710), .A2(img[504]), .B1(n19388), .B2(img[376]), .O(
        n18451) );
  AOI22S U21055 ( .A1(n13833), .A2(img[248]), .B1(n18832), .B2(img[120]), .O(
        n18450) );
  AOI22S U21056 ( .A1(n19326), .A2(img[1016]), .B1(n13797), .B2(img[888]), .O(
        n18449) );
  AOI22S U21057 ( .A1(n20032), .A2(img[760]), .B1(n19709), .B2(img[632]), .O(
        n18448) );
  AN4S U21058 ( .I1(n18451), .I2(n18450), .I3(n18449), .I4(n18448), .O(n18457)
         );
  AOI22S U21059 ( .A1(n13786), .A2(img[2040]), .B1(n13794), .B2(img[1912]), 
        .O(n18455) );
  AOI22S U21060 ( .A1(n19193), .A2(img[1784]), .B1(n13798), .B2(img[1656]), 
        .O(n18454) );
  AOI22S U21061 ( .A1(n13854), .A2(img[1528]), .B1(n19955), .B2(img[1400]), 
        .O(n18453) );
  AOI22S U21062 ( .A1(n14189), .A2(img[1272]), .B1(n13893), .B2(img[1144]), 
        .O(n18452) );
  AN4S U21063 ( .I1(n18455), .I2(n18454), .I3(n18453), .I4(n18452), .O(n18456)
         );
  AOI22S U21064 ( .A1(n19824), .A2(n13804), .B1(n13846), .B2(n20344), .O(
        n18479) );
  AOI22S U21065 ( .A1(n19342), .A2(img[984]), .B1(n13797), .B2(img[856]), .O(
        n18461) );
  AOI22S U21066 ( .A1(n19343), .A2(img[728]), .B1(n13879), .B2(img[600]), .O(
        n18460) );
  AOI22S U21067 ( .A1(n19344), .A2(img[472]), .B1(n13836), .B2(img[344]), .O(
        n18459) );
  AOI22S U21068 ( .A1(n13801), .A2(img[216]), .B1(n20193), .B2(img[88]), .O(
        n18458) );
  AN4S U21069 ( .I1(n18461), .I2(n18460), .I3(n18459), .I4(n18458), .O(n18467)
         );
  AOI22S U21070 ( .A1(n19215), .A2(img[2008]), .B1(n13832), .B2(img[1880]), 
        .O(n18465) );
  AOI22S U21071 ( .A1(n19193), .A2(img[1752]), .B1(n17862), .B2(img[1624]), 
        .O(n18464) );
  AOI22S U21072 ( .A1(n17088), .A2(img[1496]), .B1(n19349), .B2(img[1368]), 
        .O(n18463) );
  AOI22S U21073 ( .A1(n16515), .A2(img[1240]), .B1(n13893), .B2(img[1112]), 
        .O(n18462) );
  AN4S U21074 ( .I1(n18465), .I2(n18464), .I3(n18463), .I4(n18462), .O(n18466)
         );
  ND2 U21075 ( .I1(n18467), .I2(n18466), .O(n19828) );
  AOI22S U21076 ( .A1(n19326), .A2(img[992]), .B1(n13837), .B2(img[864]), .O(
        n18471) );
  AOI22S U21077 ( .A1(n19343), .A2(img[736]), .B1(n13896), .B2(img[608]), .O(
        n18470) );
  AOI22S U21078 ( .A1(n19410), .A2(img[480]), .B1(n13836), .B2(img[352]), .O(
        n18469) );
  AOI22S U21079 ( .A1(n19290), .A2(img[224]), .B1(n20193), .B2(img[96]), .O(
        n18468) );
  AN4S U21080 ( .I1(n18471), .I2(n18470), .I3(n18469), .I4(n18468), .O(n18477)
         );
  AOI22S U21081 ( .A1(n13786), .A2(img[2016]), .B1(n18201), .B2(img[1888]), 
        .O(n18475) );
  AOI22S U21082 ( .A1(n19193), .A2(img[1760]), .B1(n17862), .B2(img[1632]), 
        .O(n18474) );
  AOI22S U21083 ( .A1(n17336), .A2(img[1504]), .B1(n19417), .B2(img[1376]), 
        .O(n18473) );
  AOI22S U21084 ( .A1(n17810), .A2(img[1248]), .B1(n13890), .B2(img[1120]), 
        .O(n18472) );
  AN4S U21085 ( .I1(n18475), .I2(n18474), .I3(n18473), .I4(n18472), .O(n18476)
         );
  ND2 U21086 ( .I1(n18477), .I2(n18476), .O(n19806) );
  AOI22S U21087 ( .A1(n19828), .A2(n17938), .B1(n13835), .B2(n19806), .O(
        n18478) );
  ND2S U21088 ( .I1(n18479), .I2(n18478), .O(n18480) );
  NR2 U21089 ( .I1(n18481), .I2(n18480), .O(n18482) );
  INV1S U21090 ( .I(n19601), .O(n18486) );
  INV1S U21091 ( .I(n20344), .O(n18485) );
  INV1S U21092 ( .I(n18142), .O(n18656) );
  OAI22S U21093 ( .A1(n18486), .A2(n18485), .B1(n18656), .B2(n18484), .O(
        n18487) );
  AOI12HS U21094 ( .B1(n20344), .B2(n19600), .A1(n18487), .O(n18488) );
  OAI12HS U21095 ( .B1(n18489), .B2(n19871), .A1(n18488), .O(n18490) );
  INV1S U21096 ( .I(n19438), .O(n18493) );
  MOAI1H U21097 ( .A1(n22940), .A2(n13822), .B1(n20345), .B2(n18493), .O(
        n21649) );
  INV4 U21098 ( .I(n21649), .O(n27893) );
  AN2 U21099 ( .I1(n21809), .I2(n20809), .O(n21635) );
  ND2T U21100 ( .I1(n21810), .I2(n20809), .O(n29461) );
  AOI22S U21101 ( .A1(n19288), .A2(img[1009]), .B1(n13797), .B2(img[881]), .O(
        n18497) );
  AOI22S U21102 ( .A1(n13785), .A2(img[753]), .B1(n13858), .B2(img[625]), .O(
        n18496) );
  AOI22S U21103 ( .A1(n19710), .A2(img[497]), .B1(n19388), .B2(img[369]), .O(
        n18495) );
  AOI22S U21104 ( .A1(n18773), .A2(img[241]), .B1(n18832), .B2(img[113]), .O(
        n18494) );
  AN4S U21105 ( .I1(n18497), .I2(n18496), .I3(n18495), .I4(n18494), .O(n18503)
         );
  AOI22S U21106 ( .A1(n19215), .A2(img[2033]), .B1(n13794), .B2(img[1905]), 
        .O(n18501) );
  AOI22S U21107 ( .A1(n13823), .A2(img[1777]), .B1(n13845), .B2(img[1649]), 
        .O(n18500) );
  AOI22S U21108 ( .A1(n13783), .A2(img[1521]), .B1(n15800), .B2(img[1393]), 
        .O(n18499) );
  AOI22S U21109 ( .A1(n13788), .A2(img[1265]), .B1(n13893), .B2(img[1137]), 
        .O(n18498) );
  AOI22S U21110 ( .A1(n16348), .A2(img[945]), .B1(n13797), .B2(img[817]), .O(
        n18507) );
  AOI22S U21111 ( .A1(n20102), .A2(img[689]), .B1(n13855), .B2(img[561]), .O(
        n18506) );
  AOI22S U21112 ( .A1(n18818), .A2(img[433]), .B1(n17611), .B2(img[305]), .O(
        n18505) );
  BUF4 U21113 ( .I(n17514), .O(n18832) );
  AOI22S U21114 ( .A1(n17793), .A2(img[177]), .B1(n18832), .B2(img[49]), .O(
        n18504) );
  AN4S U21115 ( .I1(n18507), .I2(n18506), .I3(n18505), .I4(n18504), .O(n18513)
         );
  AOI22S U21116 ( .A1(n13786), .A2(img[1969]), .B1(n19715), .B2(img[1841]), 
        .O(n18511) );
  AOI22S U21117 ( .A1(n19193), .A2(img[1713]), .B1(n13799), .B2(img[1585]), 
        .O(n18510) );
  INV1S U21118 ( .I(n13789), .O(n18729) );
  AOI22S U21119 ( .A1(n18729), .A2(img[1457]), .B1(n19647), .B2(img[1329]), 
        .O(n18509) );
  AOI22S U21120 ( .A1(n18148), .A2(img[1201]), .B1(n13889), .B2(img[1073]), 
        .O(n18508) );
  AN4S U21121 ( .I1(n18511), .I2(n18510), .I3(n18509), .I4(n18508), .O(n18512)
         );
  ND2P U21122 ( .I1(n18513), .I2(n18512), .O(n19759) );
  AOI22S U21123 ( .A1(n19770), .A2(n13839), .B1(n17875), .B2(n19759), .O(
        n18578) );
  AOI22S U21124 ( .A1(n13826), .A2(img[1001]), .B1(n13837), .B2(img[873]), .O(
        n18517) );
  AOI22S U21125 ( .A1(n19343), .A2(img[745]), .B1(n13858), .B2(img[617]), .O(
        n18516) );
  BUF1 U21126 ( .I(n13800), .O(n18831) );
  AOI22S U21127 ( .A1(n18831), .A2(img[489]), .B1(n17611), .B2(img[361]), .O(
        n18515) );
  AOI22S U21128 ( .A1(n18773), .A2(img[233]), .B1(n18832), .B2(img[105]), .O(
        n18514) );
  AN4S U21129 ( .I1(n18517), .I2(n18516), .I3(n18515), .I4(n18514), .O(n18523)
         );
  AOI22S U21130 ( .A1(n19036), .A2(img[2025]), .B1(n19416), .B2(img[1897]), 
        .O(n18521) );
  AOI22S U21131 ( .A1(n18837), .A2(img[1769]), .B1(n17862), .B2(img[1641]), 
        .O(n18520) );
  AOI22S U21132 ( .A1(n13824), .A2(img[1513]), .B1(n18838), .B2(img[1385]), 
        .O(n18519) );
  AOI22S U21133 ( .A1(n17810), .A2(img[1257]), .B1(n13861), .B2(img[1129]), 
        .O(n18518) );
  AOI22S U21134 ( .A1(n18702), .A2(img[953]), .B1(n13797), .B2(img[825]), .O(
        n18527) );
  AOI22S U21135 ( .A1(n18681), .A2(img[697]), .B1(n13896), .B2(img[569]), .O(
        n18526) );
  AOI22S U21136 ( .A1(n13829), .A2(img[441]), .B1(n17611), .B2(img[313]), .O(
        n18525) );
  AOI22S U21137 ( .A1(n13803), .A2(img[185]), .B1(n18832), .B2(img[57]), .O(
        n18524) );
  AN4S U21138 ( .I1(n18527), .I2(n18526), .I3(n18525), .I4(n18524), .O(n18533)
         );
  BUF1 U21139 ( .I(n14044), .O(n19416) );
  AOI22S U21140 ( .A1(n19036), .A2(img[1977]), .B1(n19416), .B2(img[1849]), 
        .O(n18531) );
  AOI22S U21141 ( .A1(n17382), .A2(img[1721]), .B1(n18751), .B2(img[1593]), 
        .O(n18530) );
  AOI22S U21142 ( .A1(n18298), .A2(img[1465]), .B1(n17712), .B2(img[1337]), 
        .O(n18529) );
  AOI22S U21143 ( .A1(n18935), .A2(img[1209]), .B1(n13893), .B2(img[1081]), 
        .O(n18528) );
  AN4S U21144 ( .I1(n18531), .I2(n18530), .I3(n18529), .I4(n18528), .O(n18532)
         );
  AOI22S U21145 ( .A1(n19754), .A2(n19483), .B1(n20187), .B2(n19758), .O(
        n18577) );
  AOI22S U21146 ( .A1(n19342), .A2(img[961]), .B1(n13837), .B2(img[833]), .O(
        n18537) );
  AOI22S U21147 ( .A1(n20102), .A2(img[705]), .B1(n13855), .B2(img[577]), .O(
        n18536) );
  AOI22S U21148 ( .A1(n18713), .A2(img[449]), .B1(n17611), .B2(img[321]), .O(
        n18535) );
  AOI22S U21149 ( .A1(n13803), .A2(img[193]), .B1(n18832), .B2(img[65]), .O(
        n18534) );
  AN4S U21150 ( .I1(n18537), .I2(n18536), .I3(n18535), .I4(n18534), .O(n18543)
         );
  AOI22S U21151 ( .A1(n19036), .A2(img[1985]), .B1(n18201), .B2(img[1857]), 
        .O(n18541) );
  AOI22S U21152 ( .A1(n17382), .A2(img[1729]), .B1(n17862), .B2(img[1601]), 
        .O(n18540) );
  AOI22S U21153 ( .A1(n13824), .A2(img[1473]), .B1(n18548), .B2(img[1345]), 
        .O(n18539) );
  AOI22S U21154 ( .A1(n19956), .A2(img[1217]), .B1(n13890), .B2(img[1089]), 
        .O(n18538) );
  AN4S U21155 ( .I1(n18541), .I2(n18540), .I3(n18539), .I4(n18538), .O(n18542)
         );
  AOI22S U21156 ( .A1(n16348), .A2(img[937]), .B1(n13898), .B2(img[809]), .O(
        n18547) );
  AOI22S U21157 ( .A1(n18681), .A2(img[681]), .B1(n13855), .B2(img[553]), .O(
        n18546) );
  AOI22S U21158 ( .A1(n18772), .A2(img[425]), .B1(n17611), .B2(img[297]), .O(
        n18545) );
  AOI22S U21159 ( .A1(n18958), .A2(img[169]), .B1(n18832), .B2(img[41]), .O(
        n18544) );
  AN4S U21160 ( .I1(n18547), .I2(n18546), .I3(n18545), .I4(n18544), .O(n18554)
         );
  AOI22S U21161 ( .A1(n19036), .A2(img[1961]), .B1(n19416), .B2(img[1833]), 
        .O(n18552) );
  AOI22S U21162 ( .A1(n17382), .A2(img[1705]), .B1(n18751), .B2(img[1577]), 
        .O(n18551) );
  AOI22S U21163 ( .A1(n17312), .A2(img[1449]), .B1(n18548), .B2(img[1321]), 
        .O(n18550) );
  AOI22S U21164 ( .A1(n16515), .A2(img[1193]), .B1(n13877), .B2(img[1065]), 
        .O(n18549) );
  AN4S U21165 ( .I1(n18552), .I2(n18551), .I3(n18550), .I4(n18549), .O(n18553)
         );
  ND2P U21166 ( .I1(n18554), .I2(n18553), .O(n19757) );
  AOI22S U21167 ( .A1(n19756), .A2(n13843), .B1(n20124), .B2(n19757), .O(
        n18576) );
  AOI22S U21168 ( .A1(n19641), .A2(img[969]), .B1(n13797), .B2(img[841]), .O(
        n18558) );
  AOI22S U21169 ( .A1(n13876), .A2(img[713]), .B1(n13858), .B2(img[585]), .O(
        n18557) );
  BUF1 U21170 ( .I(n13800), .O(n18736) );
  AOI22S U21171 ( .A1(n18736), .A2(img[457]), .B1(n17611), .B2(img[329]), .O(
        n18556) );
  AOI22S U21172 ( .A1(n14909), .A2(img[201]), .B1(n18832), .B2(img[73]), .O(
        n18555) );
  AN4S U21173 ( .I1(n18558), .I2(n18557), .I3(n18556), .I4(n18555), .O(n18564)
         );
  AOI22S U21174 ( .A1(n19215), .A2(img[1993]), .B1(n19715), .B2(img[1865]), 
        .O(n18562) );
  AOI22S U21175 ( .A1(n17382), .A2(img[1737]), .B1(n13845), .B2(img[1609]), 
        .O(n18561) );
  INV1S U21176 ( .I(n13789), .O(n18824) );
  AOI22S U21177 ( .A1(n18824), .A2(img[1481]), .B1(n13792), .B2(img[1353]), 
        .O(n18560) );
  AOI22S U21178 ( .A1(n16515), .A2(img[1225]), .B1(n13893), .B2(img[1097]), 
        .O(n18559) );
  AN4S U21179 ( .I1(n18562), .I2(n18561), .I3(n18560), .I4(n18559), .O(n18563)
         );
  AOI22S U21180 ( .A1(n13826), .A2(img[913]), .B1(n13797), .B2(img[785]), .O(
        n18568) );
  AOI22S U21181 ( .A1(n18681), .A2(img[657]), .B1(n13858), .B2(img[529]), .O(
        n18567) );
  BUF1 U21182 ( .I(n13800), .O(n18772) );
  AOI22S U21183 ( .A1(n18772), .A2(img[401]), .B1(n17611), .B2(img[273]), .O(
        n18566) );
  AOI22S U21184 ( .A1(n17886), .A2(img[145]), .B1(n18832), .B2(img[17]), .O(
        n18565) );
  AN4S U21185 ( .I1(n18568), .I2(n18567), .I3(n18566), .I4(n18565), .O(n18574)
         );
  AOI22S U21186 ( .A1(n19036), .A2(img[1937]), .B1(n19715), .B2(img[1809]), 
        .O(n18572) );
  AOI22S U21187 ( .A1(n17382), .A2(img[1681]), .B1(n17862), .B2(img[1553]), 
        .O(n18571) );
  INV1S U21188 ( .I(n13789), .O(n18778) );
  AOI22S U21189 ( .A1(n18778), .A2(img[1425]), .B1(n17745), .B2(img[1297]), 
        .O(n18570) );
  AOI22S U21190 ( .A1(n13788), .A2(img[1169]), .B1(n13893), .B2(img[1041]), 
        .O(n18569) );
  AOI22S U21191 ( .A1(n19747), .A2(n18040), .B1(n13830), .B2(n19752), .O(
        n18575) );
  AN4S U21192 ( .I1(n18578), .I2(n18577), .I3(n18576), .I4(n18575), .O(n18655)
         );
  AOI22S U21193 ( .A1(n17730), .A2(img[977]), .B1(n13837), .B2(img[849]), .O(
        n18582) );
  AOI22S U21194 ( .A1(n15506), .A2(img[721]), .B1(n13858), .B2(img[593]), .O(
        n18581) );
  AOI22S U21195 ( .A1(n18736), .A2(img[465]), .B1(n17611), .B2(img[337]), .O(
        n18580) );
  AOI22S U21196 ( .A1(n13833), .A2(img[209]), .B1(n18832), .B2(img[81]), .O(
        n18579) );
  AN4S U21197 ( .I1(n18582), .I2(n18581), .I3(n18580), .I4(n18579), .O(n18588)
         );
  AOI22S U21198 ( .A1(n19215), .A2(img[2001]), .B1(n19416), .B2(img[1873]), 
        .O(n18586) );
  AOI22S U21199 ( .A1(n17382), .A2(img[1745]), .B1(n17862), .B2(img[1617]), 
        .O(n18585) );
  AOI22S U21200 ( .A1(n13783), .A2(img[1489]), .B1(n13792), .B2(img[1361]), 
        .O(n18584) );
  AOI22S U21201 ( .A1(n18988), .A2(img[1233]), .B1(n13890), .B2(img[1105]), 
        .O(n18583) );
  AN4S U21202 ( .I1(n18586), .I2(n18585), .I3(n18584), .I4(n18583), .O(n18587)
         );
  AOI22S U21203 ( .A1(n13826), .A2(img[905]), .B1(n13837), .B2(img[777]), .O(
        n18592) );
  AOI22S U21204 ( .A1(n15506), .A2(img[649]), .B1(n19709), .B2(img[521]), .O(
        n18591) );
  AOI22S U21205 ( .A1(n18772), .A2(img[393]), .B1(n17611), .B2(img[265]), .O(
        n18590) );
  AOI22S U21206 ( .A1(n13833), .A2(img[137]), .B1(n18832), .B2(img[9]), .O(
        n18589) );
  AN4S U21207 ( .I1(n18592), .I2(n18591), .I3(n18590), .I4(n18589), .O(n18598)
         );
  AOI22S U21208 ( .A1(n18885), .A2(img[1929]), .B1(n19416), .B2(img[1801]), 
        .O(n18596) );
  AOI22S U21209 ( .A1(n17382), .A2(img[1673]), .B1(n17862), .B2(img[1545]), 
        .O(n18595) );
  INV1S U21210 ( .I(n13789), .O(n18789) );
  AOI22S U21211 ( .A1(n18789), .A2(img[1417]), .B1(n13787), .B2(img[1289]), 
        .O(n18594) );
  AOI22S U21212 ( .A1(n19649), .A2(img[1161]), .B1(n13893), .B2(img[1033]), 
        .O(n18593) );
  AOI22S U21213 ( .A1(n19753), .A2(n20439), .B1(n13847), .B2(n19755), .O(
        n18653) );
  AOI22S U21214 ( .A1(n13826), .A2(img[921]), .B1(n13837), .B2(img[793]), .O(
        n18602) );
  AOI22S U21215 ( .A1(n13785), .A2(img[665]), .B1(n19709), .B2(img[537]), .O(
        n18601) );
  AOI22S U21216 ( .A1(n17499), .A2(img[409]), .B1(n17611), .B2(img[281]), .O(
        n18600) );
  AOI22S U21217 ( .A1(n13841), .A2(img[153]), .B1(n18832), .B2(img[25]), .O(
        n18599) );
  AN4S U21218 ( .I1(n18602), .I2(n18601), .I3(n18600), .I4(n18599), .O(n18608)
         );
  AOI22S U21219 ( .A1(n13786), .A2(img[1945]), .B1(n19416), .B2(img[1817]), 
        .O(n18606) );
  AOI22S U21220 ( .A1(n17382), .A2(img[1689]), .B1(n17862), .B2(img[1561]), 
        .O(n18605) );
  AOI22S U21221 ( .A1(n18789), .A2(img[1433]), .B1(n18922), .B2(img[1305]), 
        .O(n18604) );
  AOI22S U21222 ( .A1(n19956), .A2(img[1177]), .B1(n13893), .B2(img[1049]), 
        .O(n18603) );
  AN4S U21223 ( .I1(n18606), .I2(n18605), .I3(n18604), .I4(n18603), .O(n18607)
         );
  ND2S U21224 ( .I1(n19743), .I2(n17762), .O(n18652) );
  AOI22S U21225 ( .A1(n13784), .A2(img[929]), .B1(n13797), .B2(img[801]), .O(
        n18612) );
  AOI22S U21226 ( .A1(n18681), .A2(img[673]), .B1(n19709), .B2(img[545]), .O(
        n18611) );
  BUF1 U21227 ( .I(n13800), .O(n18796) );
  AOI22S U21228 ( .A1(n18796), .A2(img[417]), .B1(n17611), .B2(img[289]), .O(
        n18610) );
  AOI22S U21229 ( .A1(n17793), .A2(img[161]), .B1(n18832), .B2(img[33]), .O(
        n18609) );
  AN4S U21230 ( .I1(n18612), .I2(n18611), .I3(n18610), .I4(n18609), .O(n18618)
         );
  AOI22S U21231 ( .A1(n19215), .A2(img[1953]), .B1(n19715), .B2(img[1825]), 
        .O(n18616) );
  AOI22S U21232 ( .A1(n17382), .A2(img[1697]), .B1(n18751), .B2(img[1569]), 
        .O(n18615) );
  AOI22S U21233 ( .A1(n13783), .A2(img[1441]), .B1(n18922), .B2(img[1313]), 
        .O(n18614) );
  AOI22S U21234 ( .A1(n18148), .A2(img[1185]), .B1(n13893), .B2(img[1057]), 
        .O(n18613) );
  AN4S U21235 ( .I1(n18616), .I2(n18615), .I3(n18614), .I4(n18613), .O(n18617)
         );
  AOI22S U21236 ( .A1(n19710), .A2(img[505]), .B1(n19388), .B2(img[377]), .O(
        n18622) );
  AOI22S U21237 ( .A1(n13803), .A2(img[249]), .B1(n19950), .B2(img[121]), .O(
        n18621) );
  AOI22S U21238 ( .A1(n19326), .A2(img[1017]), .B1(n13797), .B2(img[889]), .O(
        n18620) );
  AOI22S U21239 ( .A1(n20032), .A2(img[761]), .B1(n13859), .B2(img[633]), .O(
        n18619) );
  AN4S U21240 ( .I1(n18622), .I2(n18621), .I3(n18620), .I4(n18619), .O(n18629)
         );
  AOI22S U21241 ( .A1(n13867), .A2(img[2041]), .B1(n19715), .B2(img[1913]), 
        .O(n18627) );
  AOI22S U21242 ( .A1(n19193), .A2(img[1785]), .B1(n13845), .B2(img[1657]), 
        .O(n18626) );
  AOI22S U21243 ( .A1(n13854), .A2(img[1529]), .B1(n18623), .B2(img[1401]), 
        .O(n18625) );
  AOI22S U21244 ( .A1(n16515), .A2(img[1273]), .B1(n13890), .B2(img[1145]), 
        .O(n18624) );
  AOI22S U21245 ( .A1(n19744), .A2(n13804), .B1(n13846), .B2(n20324), .O(
        n18651) );
  AOI22S U21246 ( .A1(n13784), .A2(img[985]), .B1(n13797), .B2(img[857]), .O(
        n18633) );
  AOI22S U21247 ( .A1(n19343), .A2(img[729]), .B1(n13858), .B2(img[601]), .O(
        n18632) );
  AOI22S U21248 ( .A1(n18818), .A2(img[473]), .B1(n17611), .B2(img[345]), .O(
        n18631) );
  AOI22S U21249 ( .A1(n13803), .A2(img[217]), .B1(n18832), .B2(img[89]), .O(
        n18630) );
  AOI22S U21250 ( .A1(n19215), .A2(img[2009]), .B1(n19715), .B2(img[1881]), 
        .O(n18637) );
  AOI22S U21251 ( .A1(n17382), .A2(img[1753]), .B1(n13845), .B2(img[1625]), 
        .O(n18636) );
  AOI22S U21252 ( .A1(n18824), .A2(img[1497]), .B1(n18922), .B2(img[1369]), 
        .O(n18635) );
  AOI22S U21253 ( .A1(n16515), .A2(img[1241]), .B1(n13893), .B2(img[1113]), 
        .O(n18634) );
  AN4S U21254 ( .I1(n18637), .I2(n18636), .I3(n18635), .I4(n18634), .O(n18638)
         );
  AOI22S U21255 ( .A1(n13826), .A2(img[993]), .B1(n13837), .B2(img[865]), .O(
        n18643) );
  AOI22S U21256 ( .A1(n13876), .A2(img[737]), .B1(n13858), .B2(img[609]), .O(
        n18642) );
  AOI22S U21257 ( .A1(n18831), .A2(img[481]), .B1(n17611), .B2(img[353]), .O(
        n18641) );
  AOI22S U21258 ( .A1(n17816), .A2(img[225]), .B1(n18832), .B2(img[97]), .O(
        n18640) );
  AN4S U21259 ( .I1(n18643), .I2(n18642), .I3(n18641), .I4(n18640), .O(n18649)
         );
  AOI22S U21260 ( .A1(n19036), .A2(img[2017]), .B1(n13794), .B2(img[1889]), 
        .O(n18647) );
  AOI22S U21261 ( .A1(n13823), .A2(img[1761]), .B1(n13798), .B2(img[1633]), 
        .O(n18646) );
  AOI22S U21262 ( .A1(n13783), .A2(img[1505]), .B1(n18838), .B2(img[1377]), 
        .O(n18645) );
  AOI22S U21263 ( .A1(n16515), .A2(img[1249]), .B1(n13889), .B2(img[1121]), 
        .O(n18644) );
  AOI22S U21264 ( .A1(n19742), .A2(n13791), .B1(n13835), .B2(n19745), .O(
        n18650) );
  AN4S U21265 ( .I1(n18653), .I2(n18652), .I3(n18651), .I4(n18650), .O(n18654)
         );
  INV1S U21266 ( .I(n18662), .O(n18665) );
  AOI22S U21267 ( .A1(n18662), .A2(n20371), .B1(n20363), .B2(n18662), .O(
        n18664) );
  ND2S U21268 ( .I1(n20324), .I2(n19600), .O(n18660) );
  NR2 U21269 ( .I1(n20969), .I2(n18656), .O(n18658) );
  INV1S U21270 ( .I(n19554), .O(n18657) );
  AOI22S U21271 ( .A1(n18658), .A2(n18657), .B1(n19601), .B2(n20324), .O(
        n18659) );
  ND2P U21272 ( .I1(n22926), .I2(n20809), .O(n18666) );
  OAI12HP U21273 ( .B1(n15985), .B2(n19438), .A1(n18666), .O(n29475) );
  OAI22S U21274 ( .A1(n29497), .A2(n29483), .B1(n29461), .B2(n29475), .O(
        n18667) );
  AOI13HS U21275 ( .B1(n27893), .B2(n21635), .B3(n18668), .A1(n18667), .O(
        n18669) );
  NR2 U21276 ( .I1(n18670), .I2(n18669), .O(n18859) );
  INV2 U21277 ( .I(n20535), .O(n21611) );
  AOI22S U21278 ( .A1(n19342), .A2(img[1012]), .B1(n13898), .B2(img[884]), .O(
        n18674) );
  AOI22S U21279 ( .A1(n15657), .A2(img[756]), .B1(n13858), .B2(img[628]), .O(
        n18673) );
  AOI22S U21280 ( .A1(n19710), .A2(img[500]), .B1(n19388), .B2(img[372]), .O(
        n18672) );
  AOI22S U21281 ( .A1(n13801), .A2(img[244]), .B1(n18832), .B2(img[116]), .O(
        n18671) );
  AN4S U21282 ( .I1(n18674), .I2(n18673), .I3(n18672), .I4(n18671), .O(n18680)
         );
  AOI22S U21283 ( .A1(n19215), .A2(img[2036]), .B1(n19416), .B2(img[1908]), 
        .O(n18678) );
  AOI22S U21284 ( .A1(n13823), .A2(img[1780]), .B1(n19182), .B2(img[1652]), 
        .O(n18677) );
  AOI22S U21285 ( .A1(n18789), .A2(img[1524]), .B1(n15800), .B2(img[1396]), 
        .O(n18676) );
  AOI22S U21286 ( .A1(n18946), .A2(img[1268]), .B1(n13861), .B2(img[1140]), 
        .O(n18675) );
  AOI22S U21287 ( .A1(n18702), .A2(img[948]), .B1(n13837), .B2(img[820]), .O(
        n18685) );
  AOI22S U21288 ( .A1(n18681), .A2(img[692]), .B1(n13855), .B2(img[564]), .O(
        n18684) );
  AOI22S U21289 ( .A1(n17523), .A2(img[436]), .B1(n17611), .B2(img[308]), .O(
        n18683) );
  AOI22S U21290 ( .A1(n20104), .A2(img[180]), .B1(n18832), .B2(img[52]), .O(
        n18682) );
  AOI22S U21291 ( .A1(n13786), .A2(img[1972]), .B1(n19715), .B2(img[1844]), 
        .O(n18689) );
  AOI22S U21292 ( .A1(n17382), .A2(img[1716]), .B1(n17827), .B2(img[1588]), 
        .O(n18688) );
  AOI22S U21293 ( .A1(n13824), .A2(img[1460]), .B1(n19295), .B2(img[1332]), 
        .O(n18687) );
  INV1S U21294 ( .I(n17522), .O(n18718) );
  AOI22S U21295 ( .A1(n14822), .A2(img[1204]), .B1(n13890), .B2(img[1076]), 
        .O(n18686) );
  AOI22S U21296 ( .A1(n20163), .A2(n13839), .B1(n17875), .B2(n20139), .O(
        n18761) );
  AOI22S U21297 ( .A1(n13826), .A2(img[1004]), .B1(n13797), .B2(img[876]), .O(
        n18695) );
  AOI22S U21298 ( .A1(n15506), .A2(img[748]), .B1(n18262), .B2(img[620]), .O(
        n18694) );
  AOI22S U21299 ( .A1(n13829), .A2(img[492]), .B1(n17611), .B2(img[364]), .O(
        n18693) );
  AOI22S U21300 ( .A1(n17778), .A2(img[236]), .B1(n18832), .B2(img[108]), .O(
        n18692) );
  AN4S U21301 ( .I1(n18695), .I2(n18694), .I3(n18693), .I4(n18692), .O(n18701)
         );
  AOI22S U21302 ( .A1(n19215), .A2(img[2028]), .B1(n13794), .B2(img[1900]), 
        .O(n18699) );
  AOI22S U21303 ( .A1(n19193), .A2(img[1772]), .B1(n17827), .B2(img[1644]), 
        .O(n18698) );
  AOI22S U21304 ( .A1(n13783), .A2(img[1516]), .B1(n15800), .B2(img[1388]), 
        .O(n18697) );
  AOI22S U21305 ( .A1(n13788), .A2(img[1260]), .B1(n13892), .B2(img[1132]), 
        .O(n18696) );
  ND2 U21306 ( .I1(n18701), .I2(n18700), .O(n20129) );
  AOI22S U21307 ( .A1(n18702), .A2(img[956]), .B1(n13837), .B2(img[828]), .O(
        n18706) );
  AOI22S U21308 ( .A1(n13876), .A2(img[700]), .B1(n13879), .B2(img[572]), .O(
        n18705) );
  AOI22S U21309 ( .A1(n18796), .A2(img[444]), .B1(n17611), .B2(img[316]), .O(
        n18704) );
  AOI22S U21310 ( .A1(n13833), .A2(img[188]), .B1(n18832), .B2(img[60]), .O(
        n18703) );
  AN4S U21311 ( .I1(n18706), .I2(n18705), .I3(n18704), .I4(n18703), .O(n18712)
         );
  AOI22S U21312 ( .A1(n13863), .A2(img[1980]), .B1(n19416), .B2(img[1852]), 
        .O(n18710) );
  AOI22S U21313 ( .A1(n17382), .A2(img[1724]), .B1(n18751), .B2(img[1596]), 
        .O(n18709) );
  AOI22S U21314 ( .A1(n18910), .A2(img[1468]), .B1(n19271), .B2(img[1340]), 
        .O(n18708) );
  AOI22S U21315 ( .A1(n13788), .A2(img[1212]), .B1(n13890), .B2(img[1084]), 
        .O(n18707) );
  AOI22S U21316 ( .A1(n20129), .A2(n19483), .B1(n20187), .B2(n20142), .O(
        n18760) );
  AOI22S U21317 ( .A1(n19376), .A2(img[964]), .B1(n13837), .B2(img[836]), .O(
        n18717) );
  AOI22S U21318 ( .A1(n20102), .A2(img[708]), .B1(n13855), .B2(img[580]), .O(
        n18716) );
  AOI22S U21319 ( .A1(n18713), .A2(img[452]), .B1(n17611), .B2(img[324]), .O(
        n18715) );
  AOI22S U21320 ( .A1(n18797), .A2(img[196]), .B1(n18832), .B2(img[68]), .O(
        n18714) );
  AN4S U21321 ( .I1(n18717), .I2(n18716), .I3(n18715), .I4(n18714), .O(n18724)
         );
  AOI22S U21322 ( .A1(n19215), .A2(img[1988]), .B1(n19715), .B2(img[1860]), 
        .O(n18722) );
  AOI22S U21323 ( .A1(n13824), .A2(img[1476]), .B1(n13792), .B2(img[1348]), 
        .O(n18720) );
  AOI22S U21324 ( .A1(n19037), .A2(img[1220]), .B1(n13890), .B2(img[1092]), 
        .O(n18719) );
  AN4S U21325 ( .I1(n18722), .I2(n18721), .I3(n18720), .I4(n18719), .O(n18723)
         );
  AOI22S U21326 ( .A1(n16348), .A2(img[940]), .B1(n13837), .B2(img[812]), .O(
        n18728) );
  AOI22S U21327 ( .A1(n20032), .A2(img[684]), .B1(n13879), .B2(img[556]), .O(
        n18727) );
  AOI22S U21328 ( .A1(n13800), .A2(img[428]), .B1(n19388), .B2(img[300]), .O(
        n18726) );
  AOI22S U21329 ( .A1(n13803), .A2(img[172]), .B1(n17383), .B2(img[44]), .O(
        n18725) );
  AN4S U21330 ( .I1(n18728), .I2(n18727), .I3(n18726), .I4(n18725), .O(n18735)
         );
  AOI22S U21331 ( .A1(n19036), .A2(img[1964]), .B1(n19715), .B2(img[1836]), 
        .O(n18733) );
  AOI22S U21332 ( .A1(n15630), .A2(img[1708]), .B1(n13799), .B2(img[1580]), 
        .O(n18732) );
  AOI22S U21333 ( .A1(n18729), .A2(img[1452]), .B1(n18922), .B2(img[1324]), 
        .O(n18731) );
  AOI22S U21334 ( .A1(n20110), .A2(img[1196]), .B1(n15653), .B2(img[1068]), 
        .O(n18730) );
  ND2 U21335 ( .I1(n18735), .I2(n18734), .O(n20123) );
  AOI22S U21336 ( .A1(n20151), .A2(n13843), .B1(n20124), .B2(n20123), .O(
        n18759) );
  AOI22S U21337 ( .A1(n16348), .A2(img[972]), .B1(n13797), .B2(img[844]), .O(
        n18740) );
  AOI22S U21338 ( .A1(n15506), .A2(img[716]), .B1(n13858), .B2(img[588]), .O(
        n18739) );
  AOI22S U21339 ( .A1(n18736), .A2(img[460]), .B1(n17611), .B2(img[332]), .O(
        n18738) );
  AOI22S U21340 ( .A1(n13803), .A2(img[204]), .B1(n18832), .B2(img[76]), .O(
        n18737) );
  AN4S U21341 ( .I1(n18740), .I2(n18739), .I3(n18738), .I4(n18737), .O(n18746)
         );
  AOI22S U21342 ( .A1(n19215), .A2(img[1996]), .B1(n19715), .B2(img[1868]), 
        .O(n18744) );
  AOI22S U21343 ( .A1(n17382), .A2(img[1740]), .B1(n17862), .B2(img[1612]), 
        .O(n18743) );
  AOI22S U21344 ( .A1(n15315), .A2(img[1484]), .B1(n13792), .B2(img[1356]), 
        .O(n18742) );
  AOI22S U21345 ( .A1(n19649), .A2(img[1228]), .B1(n13890), .B2(img[1100]), 
        .O(n18741) );
  AOI22S U21346 ( .A1(n18702), .A2(img[916]), .B1(n13898), .B2(img[788]), .O(
        n18750) );
  AOI22S U21347 ( .A1(n13785), .A2(img[660]), .B1(n13855), .B2(img[532]), .O(
        n18749) );
  AOI22S U21348 ( .A1(n17578), .A2(img[404]), .B1(n17611), .B2(img[276]), .O(
        n18748) );
  AOI22S U21349 ( .A1(n13833), .A2(img[148]), .B1(n18832), .B2(img[20]), .O(
        n18747) );
  AN4S U21350 ( .I1(n18750), .I2(n18749), .I3(n18748), .I4(n18747), .O(n18757)
         );
  AOI22S U21351 ( .A1(n19036), .A2(img[1940]), .B1(n19715), .B2(img[1812]), 
        .O(n18755) );
  AOI22S U21352 ( .A1(n17382), .A2(img[1684]), .B1(n18751), .B2(img[1556]), 
        .O(n18754) );
  AOI22S U21353 ( .A1(n18789), .A2(img[1428]), .B1(n18922), .B2(img[1300]), 
        .O(n18753) );
  AOI22S U21354 ( .A1(n18988), .A2(img[1172]), .B1(n13877), .B2(img[1044]), 
        .O(n18752) );
  AN4S U21355 ( .I1(n18755), .I2(n18754), .I3(n18753), .I4(n18752), .O(n18756)
         );
  AOI22S U21356 ( .A1(n20149), .A2(n18040), .B1(n13830), .B2(n20140), .O(
        n18758) );
  AN4S U21357 ( .I1(n18761), .I2(n18760), .I3(n18759), .I4(n18758), .O(n18850)
         );
  AOI22S U21358 ( .A1(n13784), .A2(img[980]), .B1(n13837), .B2(img[852]), .O(
        n18765) );
  AOI22S U21359 ( .A1(n13785), .A2(img[724]), .B1(n13858), .B2(img[596]), .O(
        n18764) );
  AOI22S U21360 ( .A1(n18818), .A2(img[468]), .B1(n17611), .B2(img[340]), .O(
        n18763) );
  AOI22S U21361 ( .A1(n19411), .A2(img[212]), .B1(n18832), .B2(img[84]), .O(
        n18762) );
  AOI22S U21362 ( .A1(n19036), .A2(img[2004]), .B1(n13794), .B2(img[1876]), 
        .O(n18769) );
  AOI22S U21363 ( .A1(n18837), .A2(img[1748]), .B1(n18751), .B2(img[1620]), 
        .O(n18768) );
  AOI22S U21364 ( .A1(n13783), .A2(img[1492]), .B1(n18922), .B2(img[1364]), 
        .O(n18767) );
  AOI22S U21365 ( .A1(n17810), .A2(img[1236]), .B1(n16048), .B2(img[1108]), 
        .O(n18766) );
  AOI22S U21366 ( .A1(n13826), .A2(img[908]), .B1(n13837), .B2(img[780]), .O(
        n18777) );
  AOI22S U21367 ( .A1(n13785), .A2(img[652]), .B1(n18262), .B2(img[524]), .O(
        n18776) );
  AOI22S U21368 ( .A1(n18772), .A2(img[396]), .B1(n17611), .B2(img[268]), .O(
        n18775) );
  AOI22S U21369 ( .A1(n18819), .A2(img[140]), .B1(n18832), .B2(img[12]), .O(
        n18774) );
  AN4 U21370 ( .I1(n18777), .I2(n18776), .I3(n18775), .I4(n18774), .O(n18784)
         );
  AOI22S U21371 ( .A1(n19036), .A2(img[1932]), .B1(n19715), .B2(img[1804]), 
        .O(n18782) );
  AOI22S U21372 ( .A1(n17382), .A2(img[1676]), .B1(n17862), .B2(img[1548]), 
        .O(n18781) );
  AOI22S U21373 ( .A1(n18778), .A2(img[1420]), .B1(n13787), .B2(img[1292]), 
        .O(n18780) );
  AOI22S U21374 ( .A1(n19649), .A2(img[1164]), .B1(n13893), .B2(img[1036]), 
        .O(n18779) );
  AOI22S U21375 ( .A1(n20153), .A2(n20263), .B1(n13847), .B2(n20143), .O(
        n18848) );
  AOI22S U21376 ( .A1(n19288), .A2(img[924]), .B1(n13837), .B2(img[796]), .O(
        n18788) );
  AOI22S U21377 ( .A1(n13883), .A2(img[668]), .B1(n13879), .B2(img[540]), .O(
        n18787) );
  AOI22S U21378 ( .A1(n17354), .A2(img[412]), .B1(n17611), .B2(img[284]), .O(
        n18786) );
  AOI22S U21379 ( .A1(n13803), .A2(img[156]), .B1(n18832), .B2(img[28]), .O(
        n18785) );
  AOI22S U21380 ( .A1(n19036), .A2(img[1948]), .B1(n19416), .B2(img[1820]), 
        .O(n18793) );
  AOI22S U21381 ( .A1(n17382), .A2(img[1692]), .B1(n13798), .B2(img[1564]), 
        .O(n18792) );
  AOI22S U21382 ( .A1(n18789), .A2(img[1436]), .B1(n18922), .B2(img[1308]), 
        .O(n18791) );
  AOI22S U21383 ( .A1(n13788), .A2(img[1180]), .B1(n15653), .B2(img[1052]), 
        .O(n18790) );
  ND2S U21384 ( .I1(n20152), .I2(n17762), .O(n18847) );
  AOI22S U21385 ( .A1(n19641), .A2(img[932]), .B1(n13837), .B2(img[804]), .O(
        n18801) );
  AOI22S U21386 ( .A1(n13785), .A2(img[676]), .B1(n13855), .B2(img[548]), .O(
        n18800) );
  AOI22S U21387 ( .A1(n18796), .A2(img[420]), .B1(n17611), .B2(img[292]), .O(
        n18799) );
  AOI22S U21388 ( .A1(n13803), .A2(img[164]), .B1(n18832), .B2(img[36]), .O(
        n18798) );
  AN4S U21389 ( .I1(n18801), .I2(n18800), .I3(n18799), .I4(n18798), .O(n18807)
         );
  AOI22S U21390 ( .A1(n13786), .A2(img[1956]), .B1(n19715), .B2(img[1828]), 
        .O(n18805) );
  AOI22S U21391 ( .A1(n17382), .A2(img[1700]), .B1(n18751), .B2(img[1572]), 
        .O(n18804) );
  AOI22S U21392 ( .A1(n18963), .A2(img[1444]), .B1(n18922), .B2(img[1316]), 
        .O(n18803) );
  AOI22S U21393 ( .A1(n13788), .A2(img[1188]), .B1(n16048), .B2(img[1060]), 
        .O(n18802) );
  AOI22S U21394 ( .A1(n19710), .A2(img[508]), .B1(n19388), .B2(img[380]), .O(
        n18811) );
  AOI22S U21395 ( .A1(n17816), .A2(img[252]), .B1(n18832), .B2(img[124]), .O(
        n18810) );
  AOI22S U21396 ( .A1(n16348), .A2(img[1020]), .B1(n13898), .B2(img[892]), .O(
        n18809) );
  AOI22S U21397 ( .A1(n20032), .A2(img[764]), .B1(n15691), .B2(img[636]), .O(
        n18808) );
  AN4S U21398 ( .I1(n18811), .I2(n18810), .I3(n18809), .I4(n18808), .O(n18817)
         );
  AOI22S U21399 ( .A1(n19036), .A2(img[2044]), .B1(n18201), .B2(img[1916]), 
        .O(n18815) );
  AOI22S U21400 ( .A1(n19193), .A2(img[1788]), .B1(n17827), .B2(img[1660]), 
        .O(n18814) );
  AOI22S U21401 ( .A1(n13854), .A2(img[1532]), .B1(n20039), .B2(img[1404]), 
        .O(n18813) );
  AOI22S U21402 ( .A1(n16515), .A2(img[1276]), .B1(n16048), .B2(img[1148]), 
        .O(n18812) );
  AOI22S U21403 ( .A1(n20141), .A2(n13804), .B1(n13846), .B2(n20365), .O(
        n18846) );
  AOI22S U21404 ( .A1(n13784), .A2(img[988]), .B1(n13898), .B2(img[860]), .O(
        n18823) );
  AOI22S U21405 ( .A1(n13825), .A2(img[732]), .B1(n13858), .B2(img[604]), .O(
        n18822) );
  AOI22S U21406 ( .A1(n18818), .A2(img[476]), .B1(n17611), .B2(img[348]), .O(
        n18821) );
  AOI22S U21407 ( .A1(n18819), .A2(img[220]), .B1(n18832), .B2(img[92]), .O(
        n18820) );
  AOI22S U21408 ( .A1(n19215), .A2(img[2012]), .B1(n19715), .B2(img[1884]), 
        .O(n18828) );
  AOI22S U21409 ( .A1(n17382), .A2(img[1756]), .B1(n19182), .B2(img[1628]), 
        .O(n18827) );
  AOI22S U21410 ( .A1(n18824), .A2(img[1500]), .B1(n18922), .B2(img[1372]), 
        .O(n18826) );
  AOI22S U21411 ( .A1(n14822), .A2(img[1244]), .B1(n13893), .B2(img[1116]), 
        .O(n18825) );
  AOI22S U21412 ( .A1(n13826), .A2(img[996]), .B1(n13837), .B2(img[868]), .O(
        n18836) );
  AOI22S U21413 ( .A1(n15506), .A2(img[740]), .B1(n13858), .B2(img[612]), .O(
        n18835) );
  AOI22S U21414 ( .A1(n18831), .A2(img[484]), .B1(n17611), .B2(img[356]), .O(
        n18834) );
  AOI22S U21415 ( .A1(n17778), .A2(img[228]), .B1(n18832), .B2(img[100]), .O(
        n18833) );
  AN4S U21416 ( .I1(n18836), .I2(n18835), .I3(n18834), .I4(n18833), .O(n18844)
         );
  AOI22S U21417 ( .A1(n19036), .A2(img[2020]), .B1(n17550), .B2(img[1892]), 
        .O(n18842) );
  AOI22S U21418 ( .A1(n18837), .A2(img[1764]), .B1(n17862), .B2(img[1636]), 
        .O(n18841) );
  AOI22S U21419 ( .A1(n15315), .A2(img[1508]), .B1(n18838), .B2(img[1380]), 
        .O(n18840) );
  AOI22S U21420 ( .A1(n17810), .A2(img[1252]), .B1(n13889), .B2(img[1124]), 
        .O(n18839) );
  AOI22S U21421 ( .A1(n20154), .A2(n17938), .B1(n13835), .B2(n20138), .O(
        n18845) );
  AN4S U21422 ( .I1(n18848), .I2(n18847), .I3(n18846), .I4(n18845), .O(n18849)
         );
  ND2 U21423 ( .I1(n18850), .I2(n18849), .O(n18853) );
  INV1S U21424 ( .I(n18853), .O(n18856) );
  AOI22S U21425 ( .A1(n18853), .A2(n20363), .B1(n20364), .B2(n18853), .O(
        n18855) );
  INV1S U21426 ( .I(n20365), .O(n18851) );
  MOAI1S U21427 ( .A1(n18851), .A2(n19430), .B1(n20365), .B2(n19601), .O(
        n18852) );
  AOI12HS U21428 ( .B1(n18853), .B2(n20373), .A1(n18852), .O(n18854) );
  OAI112HS U21429 ( .C1(n18856), .C2(n19542), .A1(n18855), .B1(n18854), .O(
        n22937) );
  ND2S U21430 ( .I1(n22937), .I2(n20809), .O(n18857) );
  MOAI1S U21431 ( .A1(n21611), .A2(n28527), .B1(n20503), .B2(n27266), .O(
        n18858) );
  MOAI1S U21432 ( .A1(n18859), .A2(n18858), .B1(n21611), .B2(n28527), .O(
        n19062) );
  AOI22S U21433 ( .A1(n17835), .A2(img[1013]), .B1(n13797), .B2(img[885]), .O(
        n18863) );
  AOI22S U21434 ( .A1(n20032), .A2(img[757]), .B1(n13858), .B2(img[629]), .O(
        n18862) );
  AOI22S U21435 ( .A1(n19710), .A2(img[501]), .B1(n19388), .B2(img[373]), .O(
        n18861) );
  AOI22S U21436 ( .A1(n13841), .A2(img[245]), .B1(n19950), .B2(img[117]), .O(
        n18860) );
  AN4S U21437 ( .I1(n18863), .I2(n18862), .I3(n18861), .I4(n18860), .O(n18869)
         );
  AOI22S U21438 ( .A1(n19215), .A2(img[2037]), .B1(n13832), .B2(img[1909]), 
        .O(n18867) );
  AOI22S U21439 ( .A1(n20109), .A2(img[1781]), .B1(n17862), .B2(img[1653]), 
        .O(n18866) );
  AOI22S U21440 ( .A1(n17277), .A2(img[1525]), .B1(n20039), .B2(img[1397]), 
        .O(n18865) );
  AOI22S U21441 ( .A1(n19956), .A2(img[1269]), .B1(n13890), .B2(img[1141]), 
        .O(n18864) );
  AN4S U21442 ( .I1(n18867), .I2(n18866), .I3(n18865), .I4(n18864), .O(n18868)
         );
  ND2P U21443 ( .I1(n18869), .I2(n18868), .O(n20080) );
  AOI22S U21444 ( .A1(n13875), .A2(img[949]), .B1(n13837), .B2(img[821]), .O(
        n18873) );
  AOI22S U21445 ( .A1(n13883), .A2(img[693]), .B1(n13858), .B2(img[565]), .O(
        n18872) );
  AOI22S U21446 ( .A1(n19710), .A2(img[437]), .B1(n17611), .B2(img[309]), .O(
        n18871) );
  AOI22S U21447 ( .A1(n20104), .A2(img[181]), .B1(n19950), .B2(img[53]), .O(
        n18870) );
  AOI22S U21448 ( .A1(n13874), .A2(img[1717]), .B1(n18751), .B2(img[1589]), 
        .O(n18876) );
  AOI22S U21449 ( .A1(n18923), .A2(img[1461]), .B1(n18922), .B2(img[1333]), 
        .O(n18875) );
  AOI22S U21450 ( .A1(n16515), .A2(img[1205]), .B1(n13890), .B2(img[1077]), 
        .O(n18874) );
  AN4 U21451 ( .I1(n18877), .I2(n18876), .I3(n18875), .I4(n18874), .O(n18878)
         );
  AOI22S U21452 ( .A1(n20080), .A2(n13839), .B1(n17875), .B2(n20069), .O(
        n18956) );
  AOI22S U21453 ( .A1(n19326), .A2(img[1005]), .B1(n13898), .B2(img[877]), .O(
        n18884) );
  AOI22S U21454 ( .A1(n15657), .A2(img[749]), .B1(n13896), .B2(img[621]), .O(
        n18883) );
  BUF1S U21455 ( .I(n19710), .O(n18880) );
  AOI22S U21456 ( .A1(n18880), .A2(img[493]), .B1(n17611), .B2(img[365]), .O(
        n18882) );
  AOI22S U21457 ( .A1(n17816), .A2(img[237]), .B1(n19950), .B2(img[109]), .O(
        n18881) );
  AN4S U21458 ( .I1(n18884), .I2(n18883), .I3(n18882), .I4(n18881), .O(n18891)
         );
  AOI22S U21459 ( .A1(n18885), .A2(img[2029]), .B1(n18201), .B2(img[1901]), 
        .O(n18889) );
  AOI22S U21460 ( .A1(n15630), .A2(img[1773]), .B1(n13845), .B2(img[1645]), 
        .O(n18888) );
  AOI22S U21461 ( .A1(n17088), .A2(img[1517]), .B1(n17767), .B2(img[1389]), 
        .O(n18887) );
  AOI22S U21462 ( .A1(n14189), .A2(img[1261]), .B1(n13893), .B2(img[1133]), 
        .O(n18886) );
  AN4S U21463 ( .I1(n18889), .I2(n18888), .I3(n18887), .I4(n18886), .O(n18890)
         );
  AOI22S U21464 ( .A1(n19326), .A2(img[957]), .B1(n13898), .B2(img[829]), .O(
        n18896) );
  AOI22S U21465 ( .A1(n15506), .A2(img[701]), .B1(n13858), .B2(img[573]), .O(
        n18895) );
  AOI22S U21466 ( .A1(n18892), .A2(img[445]), .B1(n17611), .B2(img[317]), .O(
        n18894) );
  AOI22S U21467 ( .A1(n17778), .A2(img[189]), .B1(n19950), .B2(img[61]), .O(
        n18893) );
  AN4 U21468 ( .I1(n18896), .I2(n18895), .I3(n18894), .I4(n18893), .O(n18903)
         );
  AOI22S U21469 ( .A1(n19036), .A2(img[1981]), .B1(n18201), .B2(img[1853]), 
        .O(n18901) );
  AOI22S U21470 ( .A1(n13823), .A2(img[1725]), .B1(n18751), .B2(img[1597]), 
        .O(n18900) );
  AOI22S U21471 ( .A1(n18897), .A2(img[1469]), .B1(n18922), .B2(img[1341]), 
        .O(n18899) );
  AOI22S U21472 ( .A1(n16515), .A2(img[1213]), .B1(n13890), .B2(img[1085]), 
        .O(n18898) );
  ND2P U21473 ( .I1(n18903), .I2(n18902), .O(n20082) );
  AOI22S U21474 ( .A1(n20072), .A2(n19483), .B1(n20187), .B2(n20082), .O(
        n18955) );
  AOI22S U21475 ( .A1(n19326), .A2(img[965]), .B1(n13898), .B2(img[837]), .O(
        n18908) );
  AOI22S U21476 ( .A1(n13785), .A2(img[709]), .B1(n13859), .B2(img[581]), .O(
        n18907) );
  AOI22S U21477 ( .A1(n18904), .A2(img[453]), .B1(n17611), .B2(img[325]), .O(
        n18906) );
  AOI22S U21478 ( .A1(n13801), .A2(img[197]), .B1(n19950), .B2(img[69]), .O(
        n18905) );
  AN4S U21479 ( .I1(n18908), .I2(n18907), .I3(n18906), .I4(n18905), .O(n18917)
         );
  AOI22S U21480 ( .A1(n19036), .A2(img[1989]), .B1(n19715), .B2(img[1861]), 
        .O(n18915) );
  AOI22S U21481 ( .A1(n13874), .A2(img[1733]), .B1(n17862), .B2(img[1605]), 
        .O(n18914) );
  AOI22S U21482 ( .A1(n18910), .A2(img[1477]), .B1(n18909), .B2(img[1349]), 
        .O(n18913) );
  AOI22S U21483 ( .A1(n18946), .A2(img[1221]), .B1(n13893), .B2(img[1093]), 
        .O(n18912) );
  AOI22S U21484 ( .A1(n13875), .A2(img[941]), .B1(n13898), .B2(img[813]), .O(
        n18921) );
  AOI22S U21485 ( .A1(n13785), .A2(img[685]), .B1(n13859), .B2(img[557]), .O(
        n18920) );
  AOI22S U21486 ( .A1(n19710), .A2(img[429]), .B1(n17611), .B2(img[301]), .O(
        n18919) );
  AOI22S U21487 ( .A1(n19290), .A2(img[173]), .B1(n19950), .B2(img[45]), .O(
        n18918) );
  AN4S U21488 ( .I1(n18921), .I2(n18920), .I3(n18919), .I4(n18918), .O(n18929)
         );
  AOI22S U21489 ( .A1(n19036), .A2(img[1965]), .B1(n18201), .B2(img[1837]), 
        .O(n18927) );
  AOI22S U21490 ( .A1(n19193), .A2(img[1709]), .B1(n17862), .B2(img[1581]), 
        .O(n18926) );
  AOI22S U21491 ( .A1(n18923), .A2(img[1453]), .B1(n18922), .B2(img[1325]), 
        .O(n18925) );
  AOI22S U21492 ( .A1(n18946), .A2(img[1197]), .B1(n13877), .B2(img[1069]), 
        .O(n18924) );
  AN4 U21493 ( .I1(n18927), .I2(n18926), .I3(n18925), .I4(n18924), .O(n18928)
         );
  AOI22S U21494 ( .A1(n20081), .A2(n13843), .B1(n20124), .B2(n20084), .O(
        n18954) );
  AOI22S U21495 ( .A1(n13875), .A2(img[973]), .B1(n13797), .B2(img[845]), .O(
        n18933) );
  AOI22S U21496 ( .A1(n13883), .A2(img[717]), .B1(n13858), .B2(img[589]), .O(
        n18932) );
  AOI22S U21497 ( .A1(n18957), .A2(img[461]), .B1(n17611), .B2(img[333]), .O(
        n18931) );
  AOI22S U21498 ( .A1(n17515), .A2(img[205]), .B1(n19950), .B2(img[77]), .O(
        n18930) );
  AN4S U21499 ( .I1(n18933), .I2(n18932), .I3(n18931), .I4(n18930), .O(n18941)
         );
  AOI22S U21500 ( .A1(n13870), .A2(img[1997]), .B1(n13794), .B2(img[1869]), 
        .O(n18939) );
  AOI22S U21501 ( .A1(n17382), .A2(img[1741]), .B1(n13845), .B2(img[1613]), 
        .O(n18938) );
  AOI22S U21502 ( .A1(n13824), .A2(img[1485]), .B1(n19349), .B2(img[1357]), 
        .O(n18937) );
  AOI22S U21503 ( .A1(n14189), .A2(img[1229]), .B1(n13893), .B2(img[1101]), 
        .O(n18936) );
  AN4S U21504 ( .I1(n18939), .I2(n18938), .I3(n18937), .I4(n18936), .O(n18940)
         );
  AOI22S U21505 ( .A1(n19326), .A2(img[917]), .B1(n13837), .B2(img[789]), .O(
        n18945) );
  AOI22S U21506 ( .A1(n18681), .A2(img[661]), .B1(n13858), .B2(img[533]), .O(
        n18944) );
  AOI22S U21507 ( .A1(n18982), .A2(img[405]), .B1(n17611), .B2(img[277]), .O(
        n18943) );
  AOI22S U21508 ( .A1(n17864), .A2(img[149]), .B1(n19950), .B2(img[21]), .O(
        n18942) );
  AN4S U21509 ( .I1(n18945), .I2(n18944), .I3(n18943), .I4(n18942), .O(n18952)
         );
  AOI22S U21510 ( .A1(n19036), .A2(img[1941]), .B1(n19416), .B2(img[1813]), 
        .O(n18950) );
  AOI22S U21511 ( .A1(n15630), .A2(img[1685]), .B1(n18751), .B2(img[1557]), 
        .O(n18949) );
  AOI22S U21512 ( .A1(n13783), .A2(img[1429]), .B1(n19271), .B2(img[1301]), 
        .O(n18948) );
  AOI22S U21513 ( .A1(n16037), .A2(img[1173]), .B1(n16048), .B2(img[1045]), 
        .O(n18947) );
  AN4S U21514 ( .I1(n18950), .I2(n18949), .I3(n18948), .I4(n18947), .O(n18951)
         );
  AOI22S U21515 ( .A1(n20083), .A2(n20968), .B1(n13830), .B2(n20075), .O(
        n18953) );
  AOI22S U21516 ( .A1(n19326), .A2(img[981]), .B1(n13837), .B2(img[853]), .O(
        n18962) );
  AOI22S U21517 ( .A1(n13825), .A2(img[725]), .B1(n13859), .B2(img[597]), .O(
        n18961) );
  AOI22S U21518 ( .A1(n18957), .A2(img[469]), .B1(n17611), .B2(img[341]), .O(
        n18960) );
  AOI22S U21519 ( .A1(n18797), .A2(img[213]), .B1(n19950), .B2(img[85]), .O(
        n18959) );
  AN4S U21520 ( .I1(n18962), .I2(n18961), .I3(n18960), .I4(n18959), .O(n18969)
         );
  AOI22S U21521 ( .A1(n19036), .A2(img[2005]), .B1(n18201), .B2(img[1877]), 
        .O(n18967) );
  AOI22S U21522 ( .A1(n13874), .A2(img[1749]), .B1(n17827), .B2(img[1621]), 
        .O(n18966) );
  AOI22S U21523 ( .A1(n18963), .A2(img[1493]), .B1(n19417), .B2(img[1365]), 
        .O(n18965) );
  AOI22S U21524 ( .A1(n18946), .A2(img[1237]), .B1(n13880), .B2(img[1109]), 
        .O(n18964) );
  AOI22S U21525 ( .A1(n19326), .A2(img[909]), .B1(n13797), .B2(img[781]), .O(
        n18973) );
  AOI22S U21526 ( .A1(n15506), .A2(img[653]), .B1(n13896), .B2(img[525]), .O(
        n18972) );
  AOI22S U21527 ( .A1(n19710), .A2(img[397]), .B1(n17611), .B2(img[269]), .O(
        n18971) );
  AOI22S U21528 ( .A1(n17515), .A2(img[141]), .B1(n19950), .B2(img[13]), .O(
        n18970) );
  AN4S U21529 ( .I1(n18973), .I2(n18972), .I3(n18971), .I4(n18970), .O(n18981)
         );
  AOI22S U21530 ( .A1(n13786), .A2(img[1933]), .B1(n19416), .B2(img[1805]), 
        .O(n18979) );
  AOI22S U21531 ( .A1(n13823), .A2(img[1677]), .B1(n17827), .B2(img[1549]), 
        .O(n18978) );
  AOI22S U21532 ( .A1(n18975), .A2(img[1421]), .B1(n18974), .B2(img[1293]), 
        .O(n18977) );
  AOI22S U21533 ( .A1(n19649), .A2(img[1165]), .B1(n13861), .B2(img[1037]), 
        .O(n18976) );
  AN4S U21534 ( .I1(n18979), .I2(n18978), .I3(n18977), .I4(n18976), .O(n18980)
         );
  AOI22S U21535 ( .A1(n20073), .A2(n20439), .B1(n13847), .B2(n20085), .O(
        n19047) );
  AOI22S U21536 ( .A1(n19326), .A2(img[925]), .B1(n13898), .B2(img[797]), .O(
        n18987) );
  AOI22S U21537 ( .A1(n13785), .A2(img[669]), .B1(n13858), .B2(img[541]), .O(
        n18986) );
  AOI22S U21538 ( .A1(n18982), .A2(img[413]), .B1(n17611), .B2(img[285]), .O(
        n18985) );
  AOI22S U21539 ( .A1(n13841), .A2(img[157]), .B1(n19950), .B2(img[29]), .O(
        n18984) );
  AN4S U21540 ( .I1(n18987), .I2(n18986), .I3(n18985), .I4(n18984), .O(n18994)
         );
  AOI22S U21541 ( .A1(n13867), .A2(img[1949]), .B1(n13796), .B2(img[1821]), 
        .O(n18992) );
  AOI22S U21542 ( .A1(n13823), .A2(img[1693]), .B1(n17862), .B2(img[1565]), 
        .O(n18991) );
  AOI22S U21543 ( .A1(n18963), .A2(img[1437]), .B1(n17767), .B2(img[1309]), 
        .O(n18990) );
  AOI22S U21544 ( .A1(n18911), .A2(img[1181]), .B1(n13861), .B2(img[1053]), 
        .O(n18989) );
  AN4S U21545 ( .I1(n18992), .I2(n18991), .I3(n18990), .I4(n18989), .O(n18993)
         );
  ND2S U21546 ( .I1(n20070), .I2(n17762), .O(n19046) );
  AOI22S U21547 ( .A1(n19326), .A2(img[933]), .B1(n13797), .B2(img[805]), .O(
        n19000) );
  AOI22S U21548 ( .A1(n13785), .A2(img[677]), .B1(n15799), .B2(img[549]), .O(
        n18999) );
  AOI22S U21549 ( .A1(n18995), .A2(img[421]), .B1(n17611), .B2(img[293]), .O(
        n18998) );
  AOI22S U21550 ( .A1(n18819), .A2(img[165]), .B1(n19950), .B2(img[37]), .O(
        n18997) );
  AN4S U21551 ( .I1(n19000), .I2(n18999), .I3(n18998), .I4(n18997), .O(n19007)
         );
  AOI22S U21552 ( .A1(n18885), .A2(img[1957]), .B1(n18201), .B2(img[1829]), 
        .O(n19005) );
  AOI22S U21553 ( .A1(n13823), .A2(img[1701]), .B1(n19001), .B2(img[1573]), 
        .O(n19004) );
  AOI22S U21554 ( .A1(n13783), .A2(img[1445]), .B1(n13792), .B2(img[1317]), 
        .O(n19003) );
  AOI22S U21555 ( .A1(n14189), .A2(img[1189]), .B1(n13893), .B2(img[1061]), 
        .O(n19002) );
  ND2P U21556 ( .I1(n19007), .I2(n19006), .O(n20087) );
  AOI22S U21557 ( .A1(n19710), .A2(img[509]), .B1(n19388), .B2(img[381]), .O(
        n19011) );
  AOI22S U21558 ( .A1(n17886), .A2(img[253]), .B1(n18832), .B2(img[125]), .O(
        n19010) );
  AOI22S U21559 ( .A1(n19326), .A2(img[1021]), .B1(n13797), .B2(img[893]), .O(
        n19009) );
  AOI22S U21560 ( .A1(n20032), .A2(img[765]), .B1(n15799), .B2(img[637]), .O(
        n19008) );
  AN4S U21561 ( .I1(n19011), .I2(n19010), .I3(n19009), .I4(n19008), .O(n19017)
         );
  AOI22S U21562 ( .A1(n13786), .A2(img[2045]), .B1(n19416), .B2(img[1917]), 
        .O(n19015) );
  AOI22S U21563 ( .A1(n13854), .A2(img[1533]), .B1(n20039), .B2(img[1405]), 
        .O(n19013) );
  AOI22S U21564 ( .A1(n13788), .A2(img[1277]), .B1(n13877), .B2(img[1149]), 
        .O(n19012) );
  AN4S U21565 ( .I1(n19015), .I2(n19014), .I3(n19013), .I4(n19012), .O(n19016)
         );
  ND2P U21566 ( .I1(n19017), .I2(n19016), .O(n20303) );
  AOI22S U21567 ( .A1(n20087), .A2(n13804), .B1(n13846), .B2(n20303), .O(
        n19045) );
  AOI22S U21568 ( .A1(n19326), .A2(img[989]), .B1(n13837), .B2(img[861]), .O(
        n19022) );
  AOI22S U21569 ( .A1(n15506), .A2(img[733]), .B1(n13858), .B2(img[605]), .O(
        n19021) );
  AOI22S U21570 ( .A1(n19018), .A2(img[477]), .B1(n17611), .B2(img[349]), .O(
        n19020) );
  AOI22S U21571 ( .A1(n17886), .A2(img[221]), .B1(n19950), .B2(img[93]), .O(
        n19019) );
  AN4S U21572 ( .I1(n19022), .I2(n19021), .I3(n19020), .I4(n19019), .O(n19030)
         );
  AOI22S U21573 ( .A1(n19023), .A2(img[2013]), .B1(n19416), .B2(img[1885]), 
        .O(n19028) );
  AOI22S U21574 ( .A1(n13874), .A2(img[1757]), .B1(n19182), .B2(img[1629]), 
        .O(n19027) );
  AOI22S U21575 ( .A1(n13824), .A2(img[1501]), .B1(n13787), .B2(img[1373]), 
        .O(n19026) );
  AOI22S U21576 ( .A1(n14505), .A2(img[1245]), .B1(n13893), .B2(img[1117]), 
        .O(n19025) );
  AOI22S U21577 ( .A1(n19326), .A2(img[997]), .B1(n13797), .B2(img[869]), .O(
        n19035) );
  AOI22S U21578 ( .A1(n13825), .A2(img[741]), .B1(n19709), .B2(img[613]), .O(
        n19034) );
  AOI22S U21579 ( .A1(n19031), .A2(img[485]), .B1(n17611), .B2(img[357]), .O(
        n19033) );
  AOI22S U21580 ( .A1(n13801), .A2(img[229]), .B1(n19950), .B2(img[101]), .O(
        n19032) );
  AN4S U21581 ( .I1(n19035), .I2(n19034), .I3(n19033), .I4(n19032), .O(n19043)
         );
  AOI22S U21582 ( .A1(n19036), .A2(img[2021]), .B1(n18201), .B2(img[1893]), 
        .O(n19041) );
  AOI22S U21583 ( .A1(n13874), .A2(img[1765]), .B1(n13845), .B2(img[1637]), 
        .O(n19040) );
  AOI22S U21584 ( .A1(n13783), .A2(img[1509]), .B1(n19955), .B2(img[1381]), 
        .O(n19039) );
  AOI22S U21585 ( .A1(n14505), .A2(img[1253]), .B1(n13893), .B2(img[1125]), 
        .O(n19038) );
  AN4S U21586 ( .I1(n19041), .I2(n19040), .I3(n19039), .I4(n19038), .O(n19042)
         );
  ND2P U21587 ( .I1(n19043), .I2(n19042), .O(n20074) );
  AOI22S U21588 ( .A1(n20086), .A2(n13791), .B1(n13835), .B2(n20074), .O(
        n19044) );
  AN4S U21589 ( .I1(n19047), .I2(n19046), .I3(n19045), .I4(n19044), .O(n19048)
         );
  ND2 U21590 ( .I1(n19049), .I2(n19048), .O(n19054) );
  INV1S U21591 ( .I(n19054), .O(n19057) );
  AOI22S U21592 ( .A1(n19054), .A2(n20371), .B1(n20364), .B2(n19054), .O(
        n19056) );
  ND2S U21593 ( .I1(n20303), .I2(n19600), .O(n19052) );
  ND2S U21594 ( .I1(n19601), .I2(n20303), .O(n19051) );
  ND3 U21595 ( .I1(n19052), .I2(n19051), .I3(n19050), .O(n19053) );
  AOI12HS U21596 ( .B1(n19054), .B2(n20373), .A1(n19053), .O(n19055) );
  OAI112HS U21597 ( .C1(n19057), .C2(n19235), .A1(n19056), .B1(n19055), .O(
        n22921) );
  BUF1 U21598 ( .I(n19059), .O(n21411) );
  OR2 U21599 ( .I1(n21595), .I2(n21411), .O(n19061) );
  AN2S U21600 ( .I1(n19059), .I2(n21595), .O(n19060) );
  AOI12HS U21601 ( .B1(n19062), .B2(n19061), .A1(n19060), .O(n19240) );
  INV1S U21602 ( .I(n21254), .O(n20950) );
  AOI22S U21603 ( .A1(n19326), .A2(img[1014]), .B1(n13837), .B2(img[886]), .O(
        n19066) );
  AOI22S U21604 ( .A1(n20102), .A2(img[758]), .B1(n13855), .B2(img[630]), .O(
        n19065) );
  AOI22S U21605 ( .A1(n19710), .A2(img[502]), .B1(n19388), .B2(img[374]), .O(
        n19064) );
  AOI22S U21606 ( .A1(n18797), .A2(img[246]), .B1(n18832), .B2(img[118]), .O(
        n19063) );
  AN4S U21607 ( .I1(n19066), .I2(n19065), .I3(n19064), .I4(n19063), .O(n19072)
         );
  AOI22S U21608 ( .A1(n13786), .A2(img[2038]), .B1(n18201), .B2(img[1910]), 
        .O(n19070) );
  AOI22S U21609 ( .A1(n17382), .A2(img[1782]), .B1(n19182), .B2(img[1654]), 
        .O(n19069) );
  AOI22S U21610 ( .A1(n16635), .A2(img[1526]), .B1(n18922), .B2(img[1398]), 
        .O(n19068) );
  AOI22S U21611 ( .A1(n13788), .A2(img[1270]), .B1(n13890), .B2(img[1142]), 
        .O(n19067) );
  AN4S U21612 ( .I1(n19070), .I2(n19069), .I3(n19068), .I4(n19067), .O(n19071)
         );
  AOI22S U21613 ( .A1(n19252), .A2(img[950]), .B1(n13898), .B2(img[822]), .O(
        n19076) );
  AOI22S U21614 ( .A1(n13785), .A2(img[694]), .B1(n13855), .B2(img[566]), .O(
        n19075) );
  AOI22S U21615 ( .A1(n19253), .A2(img[438]), .B1(n13836), .B2(img[310]), .O(
        n19074) );
  AOI22S U21616 ( .A1(n13841), .A2(img[182]), .B1(n20193), .B2(img[54]), .O(
        n19073) );
  AN4S U21617 ( .I1(n19076), .I2(n19075), .I3(n19074), .I4(n19073), .O(n19082)
         );
  AOI22S U21618 ( .A1(n13786), .A2(img[1974]), .B1(n18201), .B2(img[1846]), 
        .O(n19080) );
  AOI22S U21619 ( .A1(n17382), .A2(img[1718]), .B1(n19182), .B2(img[1590]), 
        .O(n19079) );
  AOI22S U21620 ( .A1(n16635), .A2(img[1462]), .B1(n17865), .B2(img[1334]), 
        .O(n19078) );
  AOI22S U21621 ( .A1(n13788), .A2(img[1206]), .B1(n13893), .B2(img[1078]), 
        .O(n19077) );
  AN4S U21622 ( .I1(n19080), .I2(n19079), .I3(n19078), .I4(n19077), .O(n19081)
         );
  AOI22S U21623 ( .A1(n19987), .A2(n13839), .B1(n17875), .B2(n19997), .O(
        n19147) );
  AOI22S U21624 ( .A1(n19265), .A2(img[1006]), .B1(n13797), .B2(img[878]), .O(
        n19086) );
  AOI22S U21625 ( .A1(n19343), .A2(img[750]), .B1(n19709), .B2(img[622]), .O(
        n19085) );
  AOI22S U21626 ( .A1(n19266), .A2(img[494]), .B1(n13836), .B2(img[366]), .O(
        n19084) );
  AOI22S U21627 ( .A1(n19290), .A2(img[238]), .B1(n20193), .B2(img[110]), .O(
        n19083) );
  AN4S U21628 ( .I1(n19086), .I2(n19085), .I3(n19084), .I4(n19083), .O(n19092)
         );
  AOI22S U21629 ( .A1(n13786), .A2(img[2030]), .B1(n18201), .B2(img[1902]), 
        .O(n19090) );
  AOI22S U21630 ( .A1(n17382), .A2(img[1774]), .B1(n19182), .B2(img[1646]), 
        .O(n19089) );
  AOI22S U21631 ( .A1(n17359), .A2(img[1518]), .B1(n19271), .B2(img[1390]), 
        .O(n19088) );
  AOI22S U21632 ( .A1(n20110), .A2(img[1262]), .B1(n13880), .B2(img[1134]), 
        .O(n19087) );
  AN4S U21633 ( .I1(n19090), .I2(n19089), .I3(n19088), .I4(n19087), .O(n19091)
         );
  AOI22S U21634 ( .A1(n19288), .A2(img[958]), .B1(n13797), .B2(img[830]), .O(
        n19096) );
  AOI22S U21635 ( .A1(n15657), .A2(img[702]), .B1(n19709), .B2(img[574]), .O(
        n19095) );
  AOI22S U21636 ( .A1(n19289), .A2(img[446]), .B1(n13836), .B2(img[318]), .O(
        n19094) );
  AOI22S U21637 ( .A1(n18773), .A2(img[190]), .B1(n20193), .B2(img[62]), .O(
        n19093) );
  AN4S U21638 ( .I1(n19096), .I2(n19095), .I3(n19094), .I4(n19093), .O(n19102)
         );
  AOI22S U21639 ( .A1(n19215), .A2(img[1982]), .B1(n13832), .B2(img[1854]), 
        .O(n19100) );
  AOI22S U21640 ( .A1(n17382), .A2(img[1726]), .B1(n13845), .B2(img[1598]), 
        .O(n19099) );
  AOI22S U21641 ( .A1(n13783), .A2(img[1470]), .B1(n19295), .B2(img[1342]), 
        .O(n19098) );
  AOI22S U21642 ( .A1(n19956), .A2(img[1214]), .B1(n13890), .B2(img[1086]), 
        .O(n19097) );
  AOI22S U21643 ( .A1(n19983), .A2(n19483), .B1(n20187), .B2(n19995), .O(
        n19146) );
  AOI22S U21644 ( .A1(n19288), .A2(img[966]), .B1(n13837), .B2(img[838]), .O(
        n19106) );
  AOI22S U21645 ( .A1(n18681), .A2(img[710]), .B1(n13855), .B2(img[582]), .O(
        n19105) );
  AOI22S U21646 ( .A1(n19289), .A2(img[454]), .B1(n13836), .B2(img[326]), .O(
        n19104) );
  AOI22S U21647 ( .A1(n17793), .A2(img[198]), .B1(n20193), .B2(img[70]), .O(
        n19103) );
  AN4S U21648 ( .I1(n19106), .I2(n19105), .I3(n19104), .I4(n19103), .O(n19112)
         );
  AOI22S U21649 ( .A1(n19023), .A2(img[1990]), .B1(n13832), .B2(img[1862]), 
        .O(n19110) );
  AOI22S U21650 ( .A1(n17382), .A2(img[1734]), .B1(n19182), .B2(img[1606]), 
        .O(n19109) );
  AOI22S U21651 ( .A1(n17312), .A2(img[1478]), .B1(n19295), .B2(img[1350]), 
        .O(n19108) );
  AOI22S U21652 ( .A1(n16515), .A2(img[1222]), .B1(n13893), .B2(img[1094]), 
        .O(n19107) );
  AOI22S U21653 ( .A1(n19288), .A2(img[942]), .B1(n13837), .B2(img[814]), .O(
        n19116) );
  AOI22S U21654 ( .A1(n15506), .A2(img[686]), .B1(n13855), .B2(img[558]), .O(
        n19115) );
  AOI22S U21655 ( .A1(n19302), .A2(img[430]), .B1(n13836), .B2(img[302]), .O(
        n19114) );
  AOI22S U21656 ( .A1(n17778), .A2(img[174]), .B1(n20193), .B2(img[46]), .O(
        n19113) );
  AN4S U21657 ( .I1(n19116), .I2(n19115), .I3(n19114), .I4(n19113), .O(n19122)
         );
  AOI22S U21658 ( .A1(n13786), .A2(img[1966]), .B1(n18201), .B2(img[1838]), 
        .O(n19120) );
  AOI22S U21659 ( .A1(n17382), .A2(img[1710]), .B1(n19182), .B2(img[1582]), 
        .O(n19119) );
  AOI22S U21660 ( .A1(n17254), .A2(img[1454]), .B1(n19319), .B2(img[1326]), 
        .O(n19118) );
  AOI22S U21661 ( .A1(n13788), .A2(img[1198]), .B1(n13877), .B2(img[1070]), 
        .O(n19117) );
  AN4S U21662 ( .I1(n19120), .I2(n19119), .I3(n19118), .I4(n19117), .O(n19121)
         );
  AOI22S U21663 ( .A1(n19996), .A2(n13843), .B1(n20124), .B2(n20000), .O(
        n19145) );
  AOI22S U21664 ( .A1(n19641), .A2(img[974]), .B1(n13837), .B2(img[846]), .O(
        n19126) );
  AOI22S U21665 ( .A1(n13785), .A2(img[718]), .B1(n13855), .B2(img[590]), .O(
        n19125) );
  AOI22S U21666 ( .A1(n19313), .A2(img[462]), .B1(n13836), .B2(img[334]), .O(
        n19124) );
  AOI22S U21667 ( .A1(n18996), .A2(img[206]), .B1(n20193), .B2(img[78]), .O(
        n19123) );
  AN4S U21668 ( .I1(n19126), .I2(n19125), .I3(n19124), .I4(n19123), .O(n19133)
         );
  AOI22S U21669 ( .A1(n13786), .A2(img[1998]), .B1(n18201), .B2(img[1870]), 
        .O(n19131) );
  AOI22S U21670 ( .A1(n19193), .A2(img[1742]), .B1(n19182), .B2(img[1614]), 
        .O(n19130) );
  AOI22S U21671 ( .A1(n13783), .A2(img[1486]), .B1(n19319), .B2(img[1358]), 
        .O(n19129) );
  AOI22S U21672 ( .A1(n14505), .A2(img[1230]), .B1(n13861), .B2(img[1102]), 
        .O(n19128) );
  AN4S U21673 ( .I1(n19131), .I2(n19130), .I3(n19129), .I4(n19128), .O(n19132)
         );
  AOI22S U21674 ( .A1(n19326), .A2(img[918]), .B1(n13837), .B2(img[790]), .O(
        n19137) );
  AOI22S U21675 ( .A1(n13825), .A2(img[662]), .B1(n13858), .B2(img[534]), .O(
        n19136) );
  AOI22S U21676 ( .A1(n19327), .A2(img[406]), .B1(n13836), .B2(img[278]), .O(
        n19135) );
  AOI22S U21677 ( .A1(n13841), .A2(img[150]), .B1(n20193), .B2(img[22]), .O(
        n19134) );
  AN4S U21678 ( .I1(n19137), .I2(n19136), .I3(n19135), .I4(n19134), .O(n19143)
         );
  AOI22S U21679 ( .A1(n19215), .A2(img[1942]), .B1(n17561), .B2(img[1814]), 
        .O(n19141) );
  AOI22S U21680 ( .A1(n13823), .A2(img[1686]), .B1(n18751), .B2(img[1558]), 
        .O(n19140) );
  AOI22S U21681 ( .A1(n18923), .A2(img[1430]), .B1(n13792), .B2(img[1302]), 
        .O(n19139) );
  AOI22S U21682 ( .A1(n13788), .A2(img[1174]), .B1(n13893), .B2(img[1046]), 
        .O(n19138) );
  AN4S U21683 ( .I1(n19141), .I2(n19140), .I3(n19139), .I4(n19138), .O(n19142)
         );
  ND2 U21684 ( .I1(n19143), .I2(n19142), .O(n19985) );
  AOI22S U21685 ( .A1(n19998), .A2(n20968), .B1(n13830), .B2(n19985), .O(
        n19144) );
  AN4S U21686 ( .I1(n19147), .I2(n19146), .I3(n19145), .I4(n19144), .O(n19227)
         );
  AOI22S U21687 ( .A1(n19342), .A2(img[982]), .B1(n13837), .B2(img[854]), .O(
        n19151) );
  AOI22S U21688 ( .A1(n15657), .A2(img[726]), .B1(n13879), .B2(img[598]), .O(
        n19150) );
  AOI22S U21689 ( .A1(n19344), .A2(img[470]), .B1(n13836), .B2(img[342]), .O(
        n19149) );
  AOI22S U21690 ( .A1(n13833), .A2(img[214]), .B1(n20193), .B2(img[86]), .O(
        n19148) );
  AN4S U21691 ( .I1(n19151), .I2(n19150), .I3(n19149), .I4(n19148), .O(n19157)
         );
  AOI22S U21692 ( .A1(n19215), .A2(img[2006]), .B1(n18201), .B2(img[1878]), 
        .O(n19155) );
  AOI22S U21693 ( .A1(n15630), .A2(img[1750]), .B1(n19182), .B2(img[1622]), 
        .O(n19154) );
  AOI22S U21694 ( .A1(n13783), .A2(img[1494]), .B1(n19349), .B2(img[1366]), 
        .O(n19153) );
  AOI22S U21695 ( .A1(n18148), .A2(img[1238]), .B1(n16048), .B2(img[1110]), 
        .O(n19152) );
  AN4S U21696 ( .I1(n19155), .I2(n19154), .I3(n19153), .I4(n19152), .O(n19156)
         );
  AOI22S U21697 ( .A1(n19326), .A2(img[910]), .B1(n13797), .B2(img[782]), .O(
        n19161) );
  AOI22S U21698 ( .A1(n13825), .A2(img[654]), .B1(n13855), .B2(img[526]), .O(
        n19160) );
  AOI22S U21699 ( .A1(n20192), .A2(img[398]), .B1(n13836), .B2(img[270]), .O(
        n19159) );
  AOI22S U21700 ( .A1(n18983), .A2(img[142]), .B1(n20193), .B2(img[14]), .O(
        n19158) );
  AN4S U21701 ( .I1(n19161), .I2(n19160), .I3(n19159), .I4(n19158), .O(n19167)
         );
  AOI22S U21702 ( .A1(n19215), .A2(img[1934]), .B1(n19715), .B2(img[1806]), 
        .O(n19165) );
  AOI22S U21703 ( .A1(n13874), .A2(img[1678]), .B1(n19182), .B2(img[1550]), 
        .O(n19164) );
  AOI22S U21704 ( .A1(n13783), .A2(img[1422]), .B1(n20198), .B2(img[1294]), 
        .O(n19163) );
  AOI22S U21705 ( .A1(n19037), .A2(img[1166]), .B1(n13877), .B2(img[1038]), 
        .O(n19162) );
  AN4S U21706 ( .I1(n19165), .I2(n19164), .I3(n19163), .I4(n19162), .O(n19166)
         );
  ND2 U21707 ( .I1(n19167), .I2(n19166), .O(n20001) );
  AOI22S U21708 ( .A1(n19988), .A2(n20263), .B1(n13847), .B2(n20001), .O(
        n19225) );
  AOI22S U21709 ( .A1(n19376), .A2(img[926]), .B1(n13898), .B2(img[798]), .O(
        n19171) );
  AOI22S U21710 ( .A1(n13785), .A2(img[670]), .B1(n13855), .B2(img[542]), .O(
        n19170) );
  AOI22S U21711 ( .A1(n19377), .A2(img[414]), .B1(n13836), .B2(img[286]), .O(
        n19169) );
  AOI22S U21712 ( .A1(n13833), .A2(img[158]), .B1(n20193), .B2(img[30]), .O(
        n19168) );
  AN4S U21713 ( .I1(n19171), .I2(n19170), .I3(n19169), .I4(n19168), .O(n19177)
         );
  AOI22S U21714 ( .A1(n13786), .A2(img[1950]), .B1(n18201), .B2(img[1822]), 
        .O(n19175) );
  AOI22S U21715 ( .A1(n13874), .A2(img[1694]), .B1(n13798), .B2(img[1566]), 
        .O(n19174) );
  AOI22S U21716 ( .A1(n18963), .A2(img[1438]), .B1(n13787), .B2(img[1310]), 
        .O(n19173) );
  AOI22S U21717 ( .A1(n19037), .A2(img[1182]), .B1(n13861), .B2(img[1054]), 
        .O(n19172) );
  ND2S U21718 ( .I1(n19989), .I2(n17762), .O(n19224) );
  AOI22S U21719 ( .A1(n19376), .A2(img[934]), .B1(n13837), .B2(img[806]), .O(
        n19181) );
  AOI22S U21720 ( .A1(n15657), .A2(img[678]), .B1(n13858), .B2(img[550]), .O(
        n19180) );
  AOI22S U21721 ( .A1(n19377), .A2(img[422]), .B1(n13836), .B2(img[294]), .O(
        n19179) );
  AOI22S U21722 ( .A1(n13833), .A2(img[166]), .B1(n20193), .B2(img[38]), .O(
        n19178) );
  AN4S U21723 ( .I1(n19181), .I2(n19180), .I3(n19179), .I4(n19178), .O(n19188)
         );
  AOI22S U21724 ( .A1(n13786), .A2(img[1958]), .B1(n19715), .B2(img[1830]), 
        .O(n19186) );
  AOI22S U21725 ( .A1(n15630), .A2(img[1702]), .B1(n19182), .B2(img[1574]), 
        .O(n19185) );
  AOI22S U21726 ( .A1(n17312), .A2(img[1446]), .B1(n17840), .B2(img[1318]), 
        .O(n19184) );
  AOI22S U21727 ( .A1(n16515), .A2(img[1190]), .B1(n15653), .B2(img[1062]), 
        .O(n19183) );
  AOI22S U21728 ( .A1(n19710), .A2(img[510]), .B1(n19388), .B2(img[382]), .O(
        n19192) );
  AOI22S U21729 ( .A1(n14909), .A2(img[254]), .B1(n18832), .B2(img[126]), .O(
        n19191) );
  AOI22S U21730 ( .A1(n19342), .A2(img[1022]), .B1(n13898), .B2(img[894]), .O(
        n19190) );
  AOI22S U21731 ( .A1(n20032), .A2(img[766]), .B1(n15691), .B2(img[638]), .O(
        n19189) );
  AN4S U21732 ( .I1(n19192), .I2(n19191), .I3(n19190), .I4(n19189), .O(n19199)
         );
  AOI22S U21733 ( .A1(n13863), .A2(img[2046]), .B1(n19715), .B2(img[1918]), 
        .O(n19197) );
  AOI22S U21734 ( .A1(n19193), .A2(img[1790]), .B1(n19182), .B2(img[1662]), 
        .O(n19196) );
  AOI22S U21735 ( .A1(n17088), .A2(img[1534]), .B1(n20039), .B2(img[1406]), 
        .O(n19195) );
  AOI22S U21736 ( .A1(n18988), .A2(img[1278]), .B1(n13893), .B2(img[1150]), 
        .O(n19194) );
  AN4S U21737 ( .I1(n19197), .I2(n19196), .I3(n19195), .I4(n19194), .O(n19198)
         );
  AOI22S U21738 ( .A1(n19999), .A2(n13804), .B1(n13846), .B2(n20293), .O(
        n19223) );
  AOI22S U21739 ( .A1(n19342), .A2(img[990]), .B1(n13797), .B2(img[862]), .O(
        n19204) );
  AOI22S U21740 ( .A1(n13785), .A2(img[734]), .B1(n13855), .B2(img[606]), .O(
        n19203) );
  AOI22S U21741 ( .A1(n19344), .A2(img[478]), .B1(n13836), .B2(img[350]), .O(
        n19202) );
  AOI22S U21742 ( .A1(n13841), .A2(img[222]), .B1(n20193), .B2(img[94]), .O(
        n19201) );
  AN4S U21743 ( .I1(n19204), .I2(n19203), .I3(n19202), .I4(n19201), .O(n19210)
         );
  AOI22S U21744 ( .A1(n13786), .A2(img[2014]), .B1(n18201), .B2(img[1886]), 
        .O(n19208) );
  AOI22S U21745 ( .A1(n20109), .A2(img[1758]), .B1(n17827), .B2(img[1630]), 
        .O(n19207) );
  AOI22S U21746 ( .A1(n13783), .A2(img[1502]), .B1(n19349), .B2(img[1374]), 
        .O(n19206) );
  AOI22S U21747 ( .A1(n16515), .A2(img[1246]), .B1(n13890), .B2(img[1118]), 
        .O(n19205) );
  AN4S U21748 ( .I1(n19208), .I2(n19207), .I3(n19206), .I4(n19205), .O(n19209)
         );
  AOI22S U21749 ( .A1(n19641), .A2(img[998]), .B1(n13797), .B2(img[870]), .O(
        n19214) );
  AOI22S U21750 ( .A1(n15657), .A2(img[742]), .B1(n13896), .B2(img[614]), .O(
        n19213) );
  AOI22S U21751 ( .A1(n19410), .A2(img[486]), .B1(n13836), .B2(img[358]), .O(
        n19212) );
  AOI22S U21752 ( .A1(n18983), .A2(img[230]), .B1(n20193), .B2(img[102]), .O(
        n19211) );
  AN4S U21753 ( .I1(n19214), .I2(n19213), .I3(n19212), .I4(n19211), .O(n19221)
         );
  AOI22S U21754 ( .A1(n19215), .A2(img[2022]), .B1(n18201), .B2(img[1894]), 
        .O(n19219) );
  AOI22S U21755 ( .A1(n13874), .A2(img[1766]), .B1(n19182), .B2(img[1638]), 
        .O(n19218) );
  AOI22S U21756 ( .A1(n13783), .A2(img[1510]), .B1(n19417), .B2(img[1382]), 
        .O(n19217) );
  AOI22S U21757 ( .A1(n14189), .A2(img[1254]), .B1(n13893), .B2(img[1126]), 
        .O(n19216) );
  AN4S U21758 ( .I1(n19219), .I2(n19218), .I3(n19217), .I4(n19216), .O(n19220)
         );
  ND2 U21759 ( .I1(n19221), .I2(n19220), .O(n19994) );
  AOI22S U21760 ( .A1(n19986), .A2(n17938), .B1(n13793), .B2(n19994), .O(
        n19222) );
  AN4S U21761 ( .I1(n19225), .I2(n19224), .I3(n19223), .I4(n19222), .O(n19226)
         );
  INV1S U21762 ( .I(n19232), .O(n19236) );
  AOI22S U21763 ( .A1(n19232), .A2(n20371), .B1(n20364), .B2(n19232), .O(
        n19234) );
  ND2S U21764 ( .I1(n20293), .I2(n19600), .O(n19230) );
  ND2S U21765 ( .I1(n19601), .I2(n20293), .O(n19229) );
  ND2S U21766 ( .I1(n19474), .I2(n18142), .O(n19228) );
  ND3S U21767 ( .I1(n19230), .I2(n19229), .I3(n19228), .O(n19231) );
  AOI12HS U21768 ( .B1(n19232), .B2(n20373), .A1(n19231), .O(n19233) );
  OAI112HS U21769 ( .C1(n19236), .C2(n19235), .A1(n19234), .B1(n19233), .O(
        n22919) );
  ND2S U21770 ( .I1(n22919), .I2(n20809), .O(n19237) );
  OAI12H U21771 ( .B1(n20950), .B2(n19438), .A1(n19237), .O(n21416) );
  NR2 U21772 ( .I1(n29503), .I2(n21416), .O(n19239) );
  OAI12HS U21773 ( .B1(n19240), .B2(n19239), .A1(n19238), .O(n19441) );
  INV1S U21774 ( .I(n21259), .O(n20947) );
  AOI22S U21775 ( .A1(n16348), .A2(img[1015]), .B1(n13797), .B2(img[887]), .O(
        n19244) );
  AOI22S U21776 ( .A1(n20102), .A2(img[759]), .B1(n13859), .B2(img[631]), .O(
        n19243) );
  AOI22S U21777 ( .A1(n19710), .A2(img[503]), .B1(n19388), .B2(img[375]), .O(
        n19242) );
  AOI22S U21778 ( .A1(n20104), .A2(img[247]), .B1(n18832), .B2(img[119]), .O(
        n19241) );
  AN4S U21779 ( .I1(n19244), .I2(n19243), .I3(n19242), .I4(n19241), .O(n19251)
         );
  AOI22S U21780 ( .A1(n19023), .A2(img[2039]), .B1(n13794), .B2(img[1911]), 
        .O(n19249) );
  AOI22S U21781 ( .A1(n20109), .A2(img[1783]), .B1(n16127), .B2(img[1655]), 
        .O(n19248) );
  AOI22S U21782 ( .A1(n13783), .A2(img[1527]), .B1(n20198), .B2(img[1399]), 
        .O(n19247) );
  AOI22S U21783 ( .A1(n18911), .A2(img[1271]), .B1(n13889), .B2(img[1143]), 
        .O(n19246) );
  AN4S U21784 ( .I1(n19249), .I2(n19248), .I3(n19247), .I4(n19246), .O(n19250)
         );
  AOI22S U21785 ( .A1(n19252), .A2(img[951]), .B1(n13898), .B2(img[823]), .O(
        n19257) );
  AOI22S U21786 ( .A1(n19343), .A2(img[695]), .B1(n13896), .B2(img[567]), .O(
        n19256) );
  AOI22S U21787 ( .A1(n19253), .A2(img[439]), .B1(n13836), .B2(img[311]), .O(
        n19255) );
  AOI22S U21788 ( .A1(n18996), .A2(img[183]), .B1(n20193), .B2(img[55]), .O(
        n19254) );
  AN4S U21789 ( .I1(n19257), .I2(n19256), .I3(n19255), .I4(n19254), .O(n19264)
         );
  AOI22S U21790 ( .A1(n19036), .A2(img[1975]), .B1(n13794), .B2(img[1847]), 
        .O(n19262) );
  AOI22S U21791 ( .A1(n17382), .A2(img[1719]), .B1(n16127), .B2(img[1591]), 
        .O(n19261) );
  AOI22S U21792 ( .A1(n18778), .A2(img[1463]), .B1(n17745), .B2(img[1335]), 
        .O(n19260) );
  INV1S U21793 ( .I(n17522), .O(n19258) );
  AOI22S U21794 ( .A1(n14505), .A2(img[1207]), .B1(n13880), .B2(img[1079]), 
        .O(n19259) );
  AN4S U21795 ( .I1(n19262), .I2(n19261), .I3(n19260), .I4(n19259), .O(n19263)
         );
  ND2 U21796 ( .I1(n19264), .I2(n19263), .O(n20212) );
  AOI22S U21797 ( .A1(n20244), .A2(n13839), .B1(n17875), .B2(n20212), .O(
        n19341) );
  AOI22S U21798 ( .A1(n19265), .A2(img[1007]), .B1(n13797), .B2(img[879]), .O(
        n19270) );
  AOI22S U21799 ( .A1(n15506), .A2(img[751]), .B1(n13858), .B2(img[623]), .O(
        n19269) );
  AOI22S U21800 ( .A1(n19266), .A2(img[495]), .B1(n13836), .B2(img[367]), .O(
        n19268) );
  AOI22S U21801 ( .A1(n17793), .A2(img[239]), .B1(n20193), .B2(img[111]), .O(
        n19267) );
  AN4S U21802 ( .I1(n19270), .I2(n19269), .I3(n19268), .I4(n19267), .O(n19277)
         );
  AOI22S U21803 ( .A1(n13870), .A2(img[2031]), .B1(n13794), .B2(img[1903]), 
        .O(n19275) );
  AOI22S U21804 ( .A1(n20109), .A2(img[1775]), .B1(n19182), .B2(img[1647]), 
        .O(n19274) );
  AOI22S U21805 ( .A1(n17359), .A2(img[1519]), .B1(n19271), .B2(img[1391]), 
        .O(n19273) );
  INV1S U21806 ( .I(n16516), .O(n19403) );
  AOI22S U21807 ( .A1(n16515), .A2(img[1263]), .B1(n13877), .B2(img[1135]), 
        .O(n19272) );
  AN4S U21808 ( .I1(n19275), .I2(n19274), .I3(n19273), .I4(n19272), .O(n19276)
         );
  AOI22S U21809 ( .A1(n19288), .A2(img[959]), .B1(n13837), .B2(img[831]), .O(
        n19281) );
  AOI22S U21810 ( .A1(n13876), .A2(img[703]), .B1(n13855), .B2(img[575]), .O(
        n19280) );
  AOI22S U21811 ( .A1(n19289), .A2(img[447]), .B1(n13836), .B2(img[319]), .O(
        n19279) );
  AOI22S U21812 ( .A1(n17816), .A2(img[191]), .B1(n20193), .B2(img[63]), .O(
        n19278) );
  AN4S U21813 ( .I1(n19281), .I2(n19280), .I3(n19279), .I4(n19278), .O(n19287)
         );
  AOI22S U21814 ( .A1(n13863), .A2(img[1983]), .B1(n13794), .B2(img[1855]), 
        .O(n19285) );
  AOI22S U21815 ( .A1(n17382), .A2(img[1727]), .B1(n13798), .B2(img[1599]), 
        .O(n19284) );
  AOI22S U21816 ( .A1(n18897), .A2(img[1471]), .B1(n19295), .B2(img[1343]), 
        .O(n19283) );
  AOI22S U21817 ( .A1(n18935), .A2(img[1215]), .B1(n15653), .B2(img[1087]), 
        .O(n19282) );
  AN4S U21818 ( .I1(n19285), .I2(n19284), .I3(n19283), .I4(n19282), .O(n19286)
         );
  ND2 U21819 ( .I1(n19287), .I2(n19286), .O(n20245) );
  AOI22S U21820 ( .A1(n20233), .A2(n21062), .B1(n20187), .B2(n20245), .O(
        n19340) );
  AOI22S U21821 ( .A1(n19288), .A2(img[967]), .B1(n13837), .B2(img[839]), .O(
        n19294) );
  AOI22S U21822 ( .A1(n19343), .A2(img[711]), .B1(n13855), .B2(img[583]), .O(
        n19293) );
  AOI22S U21823 ( .A1(n19289), .A2(img[455]), .B1(n13836), .B2(img[327]), .O(
        n19292) );
  AOI22S U21824 ( .A1(n18958), .A2(img[199]), .B1(n20193), .B2(img[71]), .O(
        n19291) );
  AOI22S U21825 ( .A1(n13786), .A2(img[1991]), .B1(n13794), .B2(img[1863]), 
        .O(n19299) );
  AOI22S U21826 ( .A1(n17382), .A2(img[1735]), .B1(n13799), .B2(img[1607]), 
        .O(n19298) );
  AOI22S U21827 ( .A1(n13783), .A2(img[1479]), .B1(n19295), .B2(img[1351]), 
        .O(n19297) );
  AOI22S U21828 ( .A1(n20110), .A2(img[1223]), .B1(n15653), .B2(img[1095]), 
        .O(n19296) );
  AN4S U21829 ( .I1(n19299), .I2(n19298), .I3(n19297), .I4(n19296), .O(n19300)
         );
  ND2 U21830 ( .I1(n19301), .I2(n19300), .O(n20242) );
  AOI22S U21831 ( .A1(n13785), .A2(img[687]), .B1(n13855), .B2(img[559]), .O(
        n19305) );
  AOI22S U21832 ( .A1(n19302), .A2(img[431]), .B1(n13836), .B2(img[303]), .O(
        n19304) );
  AOI22S U21833 ( .A1(n18773), .A2(img[175]), .B1(n20193), .B2(img[47]), .O(
        n19303) );
  AN4S U21834 ( .I1(n19306), .I2(n19305), .I3(n19304), .I4(n19303), .O(n19312)
         );
  AOI22S U21835 ( .A1(n20038), .A2(img[1967]), .B1(n19715), .B2(img[1839]), 
        .O(n19310) );
  AOI22S U21836 ( .A1(n17382), .A2(img[1711]), .B1(n13798), .B2(img[1583]), 
        .O(n19309) );
  AOI22S U21837 ( .A1(n18897), .A2(img[1455]), .B1(n18838), .B2(img[1327]), 
        .O(n19308) );
  AOI22S U21838 ( .A1(n19956), .A2(img[1199]), .B1(n13892), .B2(img[1071]), 
        .O(n19307) );
  AN4S U21839 ( .I1(n19310), .I2(n19309), .I3(n19308), .I4(n19307), .O(n19311)
         );
  ND2 U21840 ( .I1(n19312), .I2(n19311), .O(n20234) );
  AOI22S U21841 ( .A1(n20242), .A2(n13843), .B1(n20124), .B2(n20234), .O(
        n19339) );
  AOI22S U21842 ( .A1(n19641), .A2(img[975]), .B1(n13797), .B2(img[847]), .O(
        n19317) );
  AOI22S U21843 ( .A1(n19343), .A2(img[719]), .B1(n13855), .B2(img[591]), .O(
        n19316) );
  AOI22S U21844 ( .A1(n19313), .A2(img[463]), .B1(n13836), .B2(img[335]), .O(
        n19315) );
  AOI22S U21845 ( .A1(n18996), .A2(img[207]), .B1(n20193), .B2(img[79]), .O(
        n19314) );
  AN4S U21846 ( .I1(n19317), .I2(n19316), .I3(n19315), .I4(n19314), .O(n19325)
         );
  AOI22S U21847 ( .A1(n13865), .A2(img[1999]), .B1(n19416), .B2(img[1871]), 
        .O(n19323) );
  AOI22S U21848 ( .A1(n17382), .A2(img[1743]), .B1(n13798), .B2(img[1615]), 
        .O(n19322) );
  AOI22S U21849 ( .A1(n13783), .A2(img[1487]), .B1(n19319), .B2(img[1359]), 
        .O(n19321) );
  AOI22S U21850 ( .A1(n18946), .A2(img[1231]), .B1(n13893), .B2(img[1103]), 
        .O(n19320) );
  AN4S U21851 ( .I1(n19323), .I2(n19322), .I3(n19321), .I4(n19320), .O(n19324)
         );
  AOI22S U21852 ( .A1(n19326), .A2(img[919]), .B1(n13797), .B2(img[791]), .O(
        n19331) );
  AOI22S U21853 ( .A1(n19343), .A2(img[663]), .B1(n13858), .B2(img[535]), .O(
        n19330) );
  AOI22S U21854 ( .A1(n19327), .A2(img[407]), .B1(n13836), .B2(img[279]), .O(
        n19329) );
  AOI22S U21855 ( .A1(n19290), .A2(img[151]), .B1(n20193), .B2(img[23]), .O(
        n19328) );
  AN4S U21856 ( .I1(n19331), .I2(n19330), .I3(n19329), .I4(n19328), .O(n19337)
         );
  AOI22S U21857 ( .A1(n19036), .A2(img[1943]), .B1(n17561), .B2(img[1815]), 
        .O(n19335) );
  AOI22S U21858 ( .A1(n19193), .A2(img[1687]), .B1(n13798), .B2(img[1559]), 
        .O(n19334) );
  AOI22S U21859 ( .A1(n18824), .A2(img[1431]), .B1(n18974), .B2(img[1303]), 
        .O(n19333) );
  AOI22S U21860 ( .A1(n19037), .A2(img[1175]), .B1(n15653), .B2(img[1047]), 
        .O(n19332) );
  AN4S U21861 ( .I1(n19335), .I2(n19334), .I3(n19333), .I4(n19332), .O(n19336)
         );
  ND2 U21862 ( .I1(n19337), .I2(n19336), .O(n20229) );
  AOI22S U21863 ( .A1(n20235), .A2(n20560), .B1(n13830), .B2(n20229), .O(
        n19338) );
  AN4S U21864 ( .I1(n19341), .I2(n19340), .I3(n19339), .I4(n19338), .O(n19429)
         );
  AOI22S U21865 ( .A1(n19342), .A2(img[983]), .B1(n13837), .B2(img[855]), .O(
        n19348) );
  AOI22S U21866 ( .A1(n19343), .A2(img[727]), .B1(n13879), .B2(img[599]), .O(
        n19347) );
  AOI22S U21867 ( .A1(n19344), .A2(img[471]), .B1(n13836), .B2(img[343]), .O(
        n19346) );
  AOI22S U21868 ( .A1(n17335), .A2(img[215]), .B1(n20193), .B2(img[87]), .O(
        n19345) );
  AN4S U21869 ( .I1(n19348), .I2(n19347), .I3(n19346), .I4(n19345), .O(n19355)
         );
  AOI22S U21870 ( .A1(n19215), .A2(img[2007]), .B1(n19416), .B2(img[1879]), 
        .O(n19353) );
  AOI22S U21871 ( .A1(n20109), .A2(img[1751]), .B1(n16127), .B2(img[1623]), 
        .O(n19352) );
  AOI22S U21872 ( .A1(n13783), .A2(img[1495]), .B1(n19349), .B2(img[1367]), 
        .O(n19351) );
  AOI22S U21873 ( .A1(n17810), .A2(img[1239]), .B1(n13893), .B2(img[1111]), 
        .O(n19350) );
  AN4S U21874 ( .I1(n19353), .I2(n19352), .I3(n19351), .I4(n19350), .O(n19354)
         );
  AOI22S U21875 ( .A1(n13875), .A2(img[911]), .B1(n13797), .B2(img[783]), .O(
        n19359) );
  AOI22S U21876 ( .A1(n13785), .A2(img[655]), .B1(n13858), .B2(img[527]), .O(
        n19358) );
  AOI22S U21877 ( .A1(n20192), .A2(img[399]), .B1(n13836), .B2(img[271]), .O(
        n19357) );
  AOI22S U21878 ( .A1(n14909), .A2(img[143]), .B1(n20193), .B2(img[15]), .O(
        n19356) );
  AN4S U21879 ( .I1(n19359), .I2(n19358), .I3(n19357), .I4(n19356), .O(n19365)
         );
  AOI22S U21880 ( .A1(n13867), .A2(img[1935]), .B1(n13794), .B2(img[1807]), 
        .O(n19363) );
  AOI22S U21881 ( .A1(n15630), .A2(img[1679]), .B1(n13798), .B2(img[1551]), 
        .O(n19362) );
  AOI22S U21882 ( .A1(n18778), .A2(img[1423]), .B1(n20198), .B2(img[1295]), 
        .O(n19361) );
  AOI22S U21883 ( .A1(n17810), .A2(img[1167]), .B1(n13890), .B2(img[1039]), 
        .O(n19360) );
  AN4S U21884 ( .I1(n19363), .I2(n19362), .I3(n19361), .I4(n19360), .O(n19364)
         );
  ND2 U21885 ( .I1(n19365), .I2(n19364), .O(n20243) );
  AOI22S U21886 ( .A1(n20232), .A2(n20263), .B1(n13847), .B2(n20243), .O(
        n19427) );
  AOI22S U21887 ( .A1(n19376), .A2(img[927]), .B1(n13898), .B2(img[799]), .O(
        n19369) );
  AOI22S U21888 ( .A1(n13825), .A2(img[671]), .B1(n13858), .B2(img[543]), .O(
        n19368) );
  AOI22S U21889 ( .A1(n19377), .A2(img[415]), .B1(n13836), .B2(img[287]), .O(
        n19367) );
  AOI22S U21890 ( .A1(n13803), .A2(img[159]), .B1(n20193), .B2(img[31]), .O(
        n19366) );
  AN4S U21891 ( .I1(n19369), .I2(n19368), .I3(n19367), .I4(n19366), .O(n19375)
         );
  AOI22S U21892 ( .A1(n19215), .A2(img[1951]), .B1(n18201), .B2(img[1823]), 
        .O(n19373) );
  AOI22S U21893 ( .A1(n19193), .A2(img[1695]), .B1(n13798), .B2(img[1567]), 
        .O(n19372) );
  AOI22S U21894 ( .A1(n18923), .A2(img[1439]), .B1(n19271), .B2(img[1311]), 
        .O(n19371) );
  AOI22S U21895 ( .A1(n13788), .A2(img[1183]), .B1(n15653), .B2(img[1055]), 
        .O(n19370) );
  AN4S U21896 ( .I1(n19373), .I2(n19372), .I3(n19371), .I4(n19370), .O(n19374)
         );
  ND2 U21897 ( .I1(n19375), .I2(n19374), .O(n20231) );
  ND2S U21898 ( .I1(n20231), .I2(n17762), .O(n19426) );
  AOI22S U21899 ( .A1(n19376), .A2(img[935]), .B1(n13797), .B2(img[807]), .O(
        n19381) );
  AOI22S U21900 ( .A1(n13785), .A2(img[679]), .B1(n13858), .B2(img[551]), .O(
        n19380) );
  AOI22S U21901 ( .A1(n19377), .A2(img[423]), .B1(n13836), .B2(img[295]), .O(
        n19379) );
  AOI22S U21902 ( .A1(n13841), .A2(img[167]), .B1(n20193), .B2(img[39]), .O(
        n19378) );
  AN4S U21903 ( .I1(n19381), .I2(n19380), .I3(n19379), .I4(n19378), .O(n19387)
         );
  AOI22S U21904 ( .A1(n19215), .A2(img[1959]), .B1(n18201), .B2(img[1831]), 
        .O(n19385) );
  AOI22S U21905 ( .A1(n19193), .A2(img[1703]), .B1(n13798), .B2(img[1575]), 
        .O(n19384) );
  AOI22S U21906 ( .A1(n17336), .A2(img[1447]), .B1(n17276), .B2(img[1319]), 
        .O(n19383) );
  AOI22S U21907 ( .A1(n14189), .A2(img[1191]), .B1(n15653), .B2(img[1063]), 
        .O(n19382) );
  AN4S U21908 ( .I1(n19385), .I2(n19384), .I3(n19383), .I4(n19382), .O(n19386)
         );
  ND2 U21909 ( .I1(n19387), .I2(n19386), .O(n20241) );
  AOI22S U21910 ( .A1(n19342), .A2(img[1023]), .B1(n13797), .B2(img[895]), .O(
        n19392) );
  AOI22S U21911 ( .A1(n15506), .A2(img[767]), .B1(n19709), .B2(img[639]), .O(
        n19391) );
  AOI22S U21912 ( .A1(n19710), .A2(img[511]), .B1(n19388), .B2(img[383]), .O(
        n19390) );
  AOI22S U21913 ( .A1(n18797), .A2(img[255]), .B1(n18832), .B2(img[127]), .O(
        n19389) );
  AN4S U21914 ( .I1(n19392), .I2(n19391), .I3(n19390), .I4(n19389), .O(n19398)
         );
  AOI22S U21915 ( .A1(n19036), .A2(img[2047]), .B1(n17561), .B2(img[1919]), 
        .O(n19396) );
  AOI22S U21916 ( .A1(n19193), .A2(img[1791]), .B1(n19001), .B2(img[1663]), 
        .O(n19395) );
  AOI22S U21917 ( .A1(n16635), .A2(img[1535]), .B1(n18922), .B2(img[1407]), 
        .O(n19394) );
  AOI22S U21918 ( .A1(n19037), .A2(img[1279]), .B1(n13893), .B2(img[1151]), 
        .O(n19393) );
  ND2 U21919 ( .I1(n19398), .I2(n19397), .O(n20281) );
  AOI22S U21920 ( .A1(n20241), .A2(n13804), .B1(n13846), .B2(n20281), .O(
        n19425) );
  AOI22S U21921 ( .A1(n13784), .A2(img[991]), .B1(n13797), .B2(img[863]), .O(
        n19402) );
  AOI22S U21922 ( .A1(n13785), .A2(img[735]), .B1(n19709), .B2(img[607]), .O(
        n19401) );
  AOI22S U21923 ( .A1(n19410), .A2(img[479]), .B1(n13836), .B2(img[351]), .O(
        n19400) );
  AOI22S U21924 ( .A1(n18996), .A2(img[223]), .B1(n20193), .B2(img[95]), .O(
        n19399) );
  AN4S U21925 ( .I1(n19402), .I2(n19401), .I3(n19400), .I4(n19399), .O(n19409)
         );
  AOI22S U21926 ( .A1(n19023), .A2(img[2015]), .B1(n19715), .B2(img[1887]), 
        .O(n19407) );
  AOI22S U21927 ( .A1(n20109), .A2(img[1759]), .B1(n13798), .B2(img[1631]), 
        .O(n19406) );
  AOI22S U21928 ( .A1(n18897), .A2(img[1503]), .B1(n19417), .B2(img[1375]), 
        .O(n19405) );
  AOI22S U21929 ( .A1(n18946), .A2(img[1247]), .B1(n13877), .B2(img[1119]), 
        .O(n19404) );
  AN4S U21930 ( .I1(n19407), .I2(n19406), .I3(n19405), .I4(n19404), .O(n19408)
         );
  AOI22S U21931 ( .A1(n19265), .A2(img[999]), .B1(n13797), .B2(img[871]), .O(
        n19415) );
  AOI22S U21932 ( .A1(n15506), .A2(img[743]), .B1(n13879), .B2(img[615]), .O(
        n19414) );
  AOI22S U21933 ( .A1(n19410), .A2(img[487]), .B1(n13836), .B2(img[359]), .O(
        n19413) );
  AOI22S U21934 ( .A1(n18983), .A2(img[231]), .B1(n20193), .B2(img[103]), .O(
        n19412) );
  AOI22S U21935 ( .A1(n19036), .A2(img[2023]), .B1(n19416), .B2(img[1895]), 
        .O(n19421) );
  AOI22S U21936 ( .A1(n20109), .A2(img[1767]), .B1(n13798), .B2(img[1639]), 
        .O(n19420) );
  AOI22S U21937 ( .A1(n13783), .A2(img[1511]), .B1(n19417), .B2(img[1383]), 
        .O(n19419) );
  AOI22S U21938 ( .A1(n18988), .A2(img[1255]), .B1(n13893), .B2(img[1127]), 
        .O(n19418) );
  AN4S U21939 ( .I1(n19421), .I2(n19420), .I3(n19419), .I4(n19418), .O(n19422)
         );
  ND2S U21940 ( .I1(n19423), .I2(n19422), .O(n20211) );
  AOI22S U21941 ( .A1(n20240), .A2(n17938), .B1(n20406), .B2(n20211), .O(
        n19424) );
  AN4S U21942 ( .I1(n19427), .I2(n19426), .I3(n19425), .I4(n19424), .O(n19428)
         );
  ND2S U21943 ( .I1(n19429), .I2(n19428), .O(n19433) );
  INV1S U21944 ( .I(n19433), .O(n19436) );
  AOI22S U21945 ( .A1(n19433), .A2(n20363), .B1(n20314), .B2(n19433), .O(
        n19435) );
  INV1S U21946 ( .I(n20281), .O(n19431) );
  MOAI1S U21947 ( .A1(n19431), .A2(n19430), .B1(n20281), .B2(n19601), .O(
        n19432) );
  AOI12HS U21948 ( .B1(n19433), .B2(n20373), .A1(n19432), .O(n19434) );
  OAI112HS U21949 ( .C1(n19436), .C2(n19661), .A1(n19435), .B1(n19434), .O(
        n22915) );
  NR2 U21950 ( .I1(n21393), .I2(n21472), .O(n19624) );
  AOI22S U21951 ( .A1(n20259), .A2(n13839), .B1(n17875), .B2(n20619), .O(
        n19445) );
  AOI22S U21952 ( .A1(n20611), .A2(n19483), .B1(n20187), .B2(n20628), .O(
        n19444) );
  AOI22S U21953 ( .A1(n20606), .A2(n14257), .B1(n20124), .B2(n20610), .O(
        n19443) );
  AOI22S U21954 ( .A1(n20614), .A2(n20968), .B1(n13830), .B2(n20621), .O(
        n19442) );
  AN4S U21955 ( .I1(n19445), .I2(n19444), .I3(n19443), .I4(n19442), .O(n19451)
         );
  AOI22S U21956 ( .A1(n20607), .A2(n20263), .B1(n13847), .B2(n20624), .O(
        n19449) );
  ND2S U21957 ( .I1(n20612), .I2(n17762), .O(n19448) );
  AOI22S U21958 ( .A1(n20626), .A2(n20620), .B1(n13846), .B2(n20608), .O(
        n19447) );
  AOI22S U21959 ( .A1(n20630), .A2(n13791), .B1(n19914), .B2(n20609), .O(
        n19446) );
  INV1S U21960 ( .I(n19457), .O(n19460) );
  INV2 U21961 ( .I(n19533), .O(n19612) );
  AOI22S U21962 ( .A1(n19457), .A2(n20364), .B1(n20314), .B2(n19457), .O(
        n19459) );
  ND2S U21963 ( .I1(n20608), .I2(n19600), .O(n19455) );
  INV1S U21964 ( .I(n22923), .O(n22918) );
  AOI22S U21965 ( .A1(n19601), .A2(n21259), .B1(n20608), .B2(n22930), .O(
        n19454) );
  ND2S U21966 ( .I1(n19603), .I2(n19452), .O(n19453) );
  AOI12HS U21967 ( .B1(n19457), .B2(n19608), .A1(n19456), .O(n19458) );
  OAI112H U21968 ( .C1(n19460), .C2(n19612), .A1(n19459), .B1(n19458), .O(
        n22410) );
  INV1S U21969 ( .I(n19461), .O(n21391) );
  AOI22S U21970 ( .A1(n19929), .A2(n13839), .B1(n17875), .B2(n20569), .O(
        n19466) );
  AOI22S U21971 ( .A1(n20593), .A2(n19483), .B1(n20963), .B2(n20579), .O(
        n19465) );
  AOI22S U21972 ( .A1(n20585), .A2(n13843), .B1(n20613), .B2(n20592), .O(
        n19464) );
  AOI22S U21973 ( .A1(n20595), .A2(n20524), .B1(n13830), .B2(n20570), .O(
        n19463) );
  AN4S U21974 ( .I1(n19466), .I2(n19465), .I3(n19464), .I4(n19463), .O(n19472)
         );
  AOI22S U21975 ( .A1(n19930), .A2(n20439), .B1(n13847), .B2(n20573), .O(
        n19470) );
  ND2S U21976 ( .I1(n20594), .I2(n17762), .O(n19469) );
  AOI22S U21977 ( .A1(n20577), .A2(n13804), .B1(n13846), .B2(n19939), .O(
        n19468) );
  AOI22S U21978 ( .A1(n20581), .A2(n13791), .B1(n19914), .B2(n20588), .O(
        n19467) );
  AN4S U21979 ( .I1(n19470), .I2(n19469), .I3(n19468), .I4(n19467), .O(n19471)
         );
  ND2S U21980 ( .I1(n19472), .I2(n19471), .O(n19479) );
  INV1S U21981 ( .I(n19479), .O(n19482) );
  AOI22S U21982 ( .A1(n19479), .A2(n19533), .B1(n20314), .B2(n19479), .O(
        n19481) );
  ND2S U21983 ( .I1(n19939), .I2(n19600), .O(n19477) );
  INV2 U21984 ( .I(n29513), .O(n22920) );
  ND2S U21985 ( .I1(n19603), .I2(n19474), .O(n19475) );
  ND3 U21986 ( .I1(n19477), .I2(n19476), .I3(n19475), .O(n19478) );
  AOI12H U21987 ( .B1(n19479), .B2(n19608), .A1(n19478), .O(n19480) );
  OAI112HP U21988 ( .C1(n19482), .C2(n19661), .A1(n19481), .B1(n19480), .O(
        n22411) );
  ND2T U21989 ( .I1(n22411), .I2(n20809), .O(n29519) );
  AOI22S U21990 ( .A1(n20013), .A2(n13839), .B1(n17875), .B2(n20551), .O(
        n19487) );
  AOI22S U21991 ( .A1(n20544), .A2(n19483), .B1(n20963), .B2(n20559), .O(
        n19486) );
  AOI22S U21992 ( .A1(n20539), .A2(n13843), .B1(n20613), .B2(n20543), .O(
        n19485) );
  AOI22S U21993 ( .A1(n20546), .A2(n21061), .B1(n13830), .B2(n20552), .O(
        n19484) );
  AN4S U21994 ( .I1(n19487), .I2(n19486), .I3(n19485), .I4(n19484), .O(n19493)
         );
  AOI22S U21995 ( .A1(n20540), .A2(n20263), .B1(n13847), .B2(n20555), .O(
        n19491) );
  ND2S U21996 ( .I1(n20545), .I2(n17762), .O(n19490) );
  AOI22S U21997 ( .A1(n20557), .A2(n13804), .B1(n13846), .B2(n20541), .O(
        n19489) );
  AOI22S U21998 ( .A1(n20561), .A2(n13791), .B1(n19914), .B2(n20542), .O(
        n19488) );
  AN4S U21999 ( .I1(n19491), .I2(n19490), .I3(n19489), .I4(n19488), .O(n19492)
         );
  ND2S U22000 ( .I1(n19493), .I2(n19492), .O(n19500) );
  INV1S U22001 ( .I(n19500), .O(n19503) );
  ND2S U22002 ( .I1(n20541), .I2(n19600), .O(n19498) );
  ND2P U22003 ( .I1(n21245), .I2(n20809), .O(n19494) );
  AOI22S U22004 ( .A1(n20366), .A2(n22922), .B1(n20541), .B2(n22930), .O(
        n19497) );
  ND2S U22005 ( .I1(n19603), .I2(n19495), .O(n19496) );
  ND3 U22006 ( .I1(n19498), .I2(n19497), .I3(n19496), .O(n19499) );
  AOI12H U22007 ( .B1(n19500), .B2(n19608), .A1(n19499), .O(n19501) );
  ND2P U22008 ( .I1(n22412), .I2(n20809), .O(n20903) );
  OAI22S U22009 ( .A1(n21804), .A2(n29519), .B1(n20903), .B2(n21805), .O(
        n19621) );
  INV1S U22010 ( .I(n21595), .O(n19619) );
  AOI22S U22011 ( .A1(n19625), .A2(n13839), .B1(n17875), .B2(n20422), .O(
        n19507) );
  AOI22S U22012 ( .A1(n20412), .A2(n19483), .B1(n20963), .B2(n20418), .O(
        n19506) );
  AOI22S U22013 ( .A1(n20403), .A2(n13843), .B1(n20124), .B2(n20413), .O(
        n19505) );
  AOI22S U22014 ( .A1(n20414), .A2(n20524), .B1(n13830), .B2(n20404), .O(
        n19504) );
  AN4S U22015 ( .I1(n19507), .I2(n19506), .I3(n19505), .I4(n19504), .O(n19513)
         );
  AOI22S U22016 ( .A1(n20407), .A2(n20263), .B1(n13847), .B2(n20419), .O(
        n19511) );
  ND2S U22017 ( .I1(n20426), .I2(n17762), .O(n19510) );
  AOI22S U22018 ( .A1(n20427), .A2(n20620), .B1(n13846), .B2(n19634), .O(
        n19509) );
  AOI22S U22019 ( .A1(n20429), .A2(n13791), .B1(n19914), .B2(n20411), .O(
        n19508) );
  AN4S U22020 ( .I1(n19511), .I2(n19510), .I3(n19509), .I4(n19508), .O(n19512)
         );
  INV1S U22021 ( .I(n19519), .O(n19522) );
  AOI22S U22022 ( .A1(n19519), .A2(n20364), .B1(n20314), .B2(n19519), .O(
        n19521) );
  ND2S U22023 ( .I1(n19634), .I2(n19600), .O(n19517) );
  ND2S U22024 ( .I1(n19603), .I2(n19514), .O(n19515) );
  ND3 U22025 ( .I1(n19517), .I2(n19516), .I3(n19515), .O(n19518) );
  AOI12HS U22026 ( .B1(n19519), .B2(n19608), .A1(n19518), .O(n19520) );
  OAI112HP U22027 ( .C1(n19522), .C2(n19612), .A1(n19521), .B1(n19520), .O(
        n22415) );
  AOI22S U22028 ( .A1(n20484), .A2(n13839), .B1(n17875), .B2(n20480), .O(
        n19526) );
  AOI22S U22029 ( .A1(n20475), .A2(n19483), .B1(n20963), .B2(n20491), .O(
        n19525) );
  AOI22S U22030 ( .A1(n20468), .A2(n13843), .B1(n20124), .B2(n20474), .O(
        n19524) );
  AOI22S U22031 ( .A1(n20476), .A2(n20524), .B1(n13830), .B2(n20481), .O(
        n19523) );
  AN4S U22032 ( .I1(n19526), .I2(n19525), .I3(n19524), .I4(n19523), .O(n19532)
         );
  AOI22S U22033 ( .A1(n20469), .A2(n20263), .B1(n13847), .B2(n20485), .O(
        n19530) );
  ND2S U22034 ( .I1(n20477), .I2(n17762), .O(n19529) );
  AOI22S U22035 ( .A1(n20489), .A2(n13804), .B1(n13846), .B2(n20470), .O(
        n19528) );
  AOI22S U22036 ( .A1(n20492), .A2(n13791), .B1(n19914), .B2(n20471), .O(
        n19527) );
  AN4S U22037 ( .I1(n19530), .I2(n19529), .I3(n19528), .I4(n19527), .O(n19531)
         );
  INV1S U22038 ( .I(n19539), .O(n19543) );
  AOI22S U22039 ( .A1(n19539), .A2(n20364), .B1(n19533), .B2(n19539), .O(
        n19541) );
  ND2S U22040 ( .I1(n20470), .I2(n19600), .O(n19537) );
  ND2S U22041 ( .I1(n19603), .I2(n19534), .O(n19535) );
  ND3 U22042 ( .I1(n19537), .I2(n19536), .I3(n19535), .O(n19538) );
  OAI112HP U22043 ( .C1(n19543), .C2(n19542), .A1(n19541), .B1(n19540), .O(
        n22416) );
  NR2 U22044 ( .I1(n22416), .I2(n29483), .O(n19589) );
  ND2T U22045 ( .I1(n22416), .I2(n20809), .O(n20891) );
  INV1S U22046 ( .I(n20891), .O(n29492) );
  AOI22S U22047 ( .A1(n20458), .A2(n13839), .B1(n17875), .B2(n20457), .O(
        n19547) );
  AOI22S U22048 ( .A1(n20444), .A2(n19483), .B1(n20963), .B2(n20455), .O(
        n19546) );
  AOI22S U22049 ( .A1(n20440), .A2(n13843), .B1(n20613), .B2(n20445), .O(
        n19545) );
  AOI22S U22050 ( .A1(n20446), .A2(n20560), .B1(n13830), .B2(n20437), .O(
        n19544) );
  AN4S U22051 ( .I1(n19547), .I2(n19546), .I3(n19545), .I4(n19544), .O(n19553)
         );
  AOI22S U22052 ( .A1(n20442), .A2(n20439), .B1(n13847), .B2(n20456), .O(
        n19551) );
  ND2S U22053 ( .I1(n20452), .I2(n17762), .O(n19550) );
  AOI22S U22054 ( .A1(n20451), .A2(n20620), .B1(n13846), .B2(n20441), .O(
        n19549) );
  AOI22S U22055 ( .A1(n20454), .A2(n13791), .B1(n19914), .B2(n20443), .O(
        n19548) );
  AN4S U22056 ( .I1(n19551), .I2(n19550), .I3(n19549), .I4(n19548), .O(n19552)
         );
  ND2P U22057 ( .I1(n19553), .I2(n19552), .O(n19559) );
  INV1S U22058 ( .I(n19559), .O(n19562) );
  AOI22S U22059 ( .A1(n19559), .A2(n20371), .B1(n20364), .B2(n19559), .O(
        n19561) );
  ND2S U22060 ( .I1(n20441), .I2(n19600), .O(n19557) );
  ND2S U22061 ( .I1(n19603), .I2(n13844), .O(n19574) );
  ND3 U22062 ( .I1(n19557), .I2(n19556), .I3(n19555), .O(n19558) );
  AOI12H U22063 ( .B1(n19559), .B2(n19608), .A1(n19558), .O(n19560) );
  OAI112HP U22064 ( .C1(n19562), .C2(n19612), .A1(n19561), .B1(n19560), .O(
        n22417) );
  ND2S U22065 ( .I1(n29461), .I2(n22417), .O(n19584) );
  AOI22S U22066 ( .A1(n21053), .A2(n13839), .B1(n17875), .B2(n21049), .O(
        n19566) );
  AOI22S U22067 ( .A1(n21044), .A2(n19483), .B1(n20963), .B2(n21060), .O(
        n19565) );
  AOI22S U22068 ( .A1(n21037), .A2(n13843), .B1(n20613), .B2(n21043), .O(
        n19564) );
  AOI22S U22069 ( .A1(n21045), .A2(n21061), .B1(n13830), .B2(n21050), .O(
        n19563) );
  AN4S U22070 ( .I1(n19566), .I2(n19565), .I3(n19564), .I4(n19563), .O(n19572)
         );
  AOI22S U22071 ( .A1(n21038), .A2(n20263), .B1(n13847), .B2(n21054), .O(
        n19570) );
  ND2S U22072 ( .I1(n21046), .I2(n17762), .O(n19569) );
  AOI22S U22073 ( .A1(n21058), .A2(n13804), .B1(n13846), .B2(n21039), .O(
        n19568) );
  AOI22S U22074 ( .A1(n21063), .A2(n13791), .B1(n19914), .B2(n21040), .O(
        n19567) );
  AN4S U22075 ( .I1(n19570), .I2(n19569), .I3(n19568), .I4(n19567), .O(n19571)
         );
  INV1S U22076 ( .I(n19580), .O(n19583) );
  AOI22S U22077 ( .A1(n19580), .A2(n20364), .B1(n20314), .B2(n19580), .O(
        n19582) );
  ND2S U22078 ( .I1(n21039), .I2(n19600), .O(n19578) );
  AOI22S U22079 ( .A1(n19601), .A2(n19573), .B1(n21039), .B2(n22930), .O(
        n19577) );
  ND3S U22080 ( .I1(n19578), .I2(n19577), .I3(n19576), .O(n19579) );
  AOI12HS U22081 ( .B1(n19580), .B2(n19608), .A1(n19579), .O(n19581) );
  OAI112HP U22082 ( .C1(n19583), .C2(n19612), .A1(n19582), .B1(n19581), .O(
        n22419) );
  INV1S U22083 ( .I(n22419), .O(n20873) );
  ND3S U22084 ( .I1(n19584), .I2(n20873), .I3(n21635), .O(n19587) );
  INV2 U22085 ( .I(n29461), .O(n20643) );
  INV1S U22086 ( .I(n22417), .O(n19585) );
  ND2S U22087 ( .I1(n20643), .I2(n19585), .O(n19586) );
  ND2T U22088 ( .I1(n22415), .I2(n20809), .O(n20892) );
  OAI22S U22089 ( .A1(n19589), .A2(n19588), .B1(n21811), .B2(n20892), .O(
        n19616) );
  AOI22S U22090 ( .A1(n20527), .A2(n13839), .B1(n17875), .B2(n20526), .O(
        n19593) );
  AOI22S U22091 ( .A1(n20512), .A2(n19483), .B1(n20963), .B2(n20523), .O(
        n19592) );
  AOI22S U22092 ( .A1(n20508), .A2(n13843), .B1(n20613), .B2(n20513), .O(
        n19591) );
  AOI22S U22093 ( .A1(n20514), .A2(n20524), .B1(n13830), .B2(n20507), .O(
        n19590) );
  AN4S U22094 ( .I1(n19593), .I2(n19592), .I3(n19591), .I4(n19590), .O(n19599)
         );
  AOI22S U22095 ( .A1(n20510), .A2(n20263), .B1(n13847), .B2(n20525), .O(
        n19597) );
  ND2S U22096 ( .I1(n20520), .I2(n17762), .O(n19596) );
  AOI22S U22097 ( .A1(n20519), .A2(n13804), .B1(n13846), .B2(n20509), .O(
        n19595) );
  AOI22S U22098 ( .A1(n20522), .A2(n13791), .B1(n19914), .B2(n20511), .O(
        n19594) );
  AN4S U22099 ( .I1(n19597), .I2(n19596), .I3(n19595), .I4(n19594), .O(n19598)
         );
  ND2S U22100 ( .I1(n19599), .I2(n19598), .O(n19609) );
  INV1S U22101 ( .I(n19609), .O(n19613) );
  AOI22S U22102 ( .A1(n19609), .A2(n20371), .B1(n20364), .B2(n19609), .O(
        n19611) );
  ND2S U22103 ( .I1(n20509), .I2(n19600), .O(n19606) );
  AOI22S U22104 ( .A1(n19601), .A2(n20863), .B1(n20509), .B2(n22930), .O(
        n19605) );
  ND2S U22105 ( .I1(n19603), .I2(n19602), .O(n19604) );
  ND3S U22106 ( .I1(n19606), .I2(n19605), .I3(n19604), .O(n19607) );
  AOI12HS U22107 ( .B1(n19609), .B2(n19608), .A1(n19607), .O(n19610) );
  OAI112H U22108 ( .C1(n19613), .C2(n19612), .A1(n19611), .B1(n19610), .O(
        n22418) );
  INV1S U22109 ( .I(n22418), .O(n19614) );
  ND2S U22110 ( .I1(n20535), .I2(n19614), .O(n19615) );
  OAI112HS U22111 ( .C1(n22415), .C2(n29442), .A1(n19616), .B1(n19615), .O(
        n19618) );
  ND2P U22112 ( .I1(n22418), .I2(n20809), .O(n20899) );
  AOI22S U22113 ( .A1(n19619), .A2(n22528), .B1(n19618), .B2(n19617), .O(
        n19620) );
  OAI22S U22114 ( .A1(n19621), .A2(n19620), .B1(n29503), .B2(n22411), .O(
        n19622) );
  OAI12HS U22115 ( .B1(n19461), .B2(n21803), .A1(n19622), .O(n19623) );
  OAI12H U22116 ( .B1(n21391), .B2(n21467), .A1(n19623), .O(n20872) );
  MOAI1 U22117 ( .A1(n19624), .A2(n20872), .B1(n21472), .B2(n21393), .O(n20662) );
  INV1S U22118 ( .I(n19625), .O(n20423) );
  MOAI1S U22119 ( .A1(n13947), .A2(n20423), .B1(n20422), .B2(n20963), .O(
        n19628) );
  INV1S U22120 ( .I(n20407), .O(n19626) );
  MOAI1S U22121 ( .A1(n13927), .A2(n19626), .B1(n20427), .B2(n20613), .O(
        n19627) );
  NR2 U22122 ( .I1(n19628), .I2(n19627), .O(n19631) );
  AOI22S U22123 ( .A1(n20414), .A2(n20439), .B1(n13793), .B2(n20429), .O(
        n19630) );
  AOI22S U22124 ( .A1(n20428), .A2(n13847), .B1(n13839), .B2(n20412), .O(
        n19629) );
  ND3S U22125 ( .I1(n19631), .I2(n19630), .I3(n19629), .O(n19708) );
  ND2S U22126 ( .I1(n20418), .I2(n17928), .O(n19633) );
  ND2S U22127 ( .I1(n20426), .I2(n20620), .O(n19632) );
  ND3S U22128 ( .I1(n19633), .I2(n19632), .I3(n13822), .O(n19636) );
  INV1S U22129 ( .I(n19634), .O(n20408) );
  MOAI1S U22130 ( .A1(n13844), .A2(n20408), .B1(n20404), .B2(n17762), .O(
        n19635) );
  NR2 U22131 ( .I1(n19636), .I2(n19635), .O(n19639) );
  AOI22S U22132 ( .A1(n20413), .A2(n17875), .B1(n13830), .B2(n20419), .O(
        n19638) );
  AOI22S U22133 ( .A1(n20411), .A2(n19483), .B1(n18040), .B2(n20403), .O(
        n19637) );
  ND3S U22134 ( .I1(n19639), .I2(n19638), .I3(n19637), .O(n19707) );
  AOI22S U22135 ( .A1(n19684), .A2(n13839), .B1(n17875), .B2(n19685), .O(
        n19640) );
  INV2 U22136 ( .I(n15142), .O(n20963) );
  AOI22S U22137 ( .A1(n19662), .A2(n20613), .B1(n17762), .B2(n19675), .O(
        n19690) );
  AOI22S U22138 ( .A1(n19665), .A2(n13830), .B1(n17928), .B2(n19674), .O(
        n19689) );
  AN4S U22139 ( .I1(n19640), .I2(n19688), .I3(n19690), .I4(n19689), .O(n19660)
         );
  AOI22S U22140 ( .A1(n19641), .A2(img[899]), .B1(n13837), .B2(img[771]), .O(
        n19646) );
  AOI22S U22141 ( .A1(n20032), .A2(img[643]), .B1(n19709), .B2(img[515]), .O(
        n19645) );
  AOI22S U22142 ( .A1(n13800), .A2(img[387]), .B1(n19388), .B2(img[259]), .O(
        n19644) );
  BUF1 U22143 ( .I(n22928), .O(n20033) );
  AOI22S U22144 ( .A1(n13833), .A2(img[131]), .B1(n20033), .B2(img[3]), .O(
        n19643) );
  AN4S U22145 ( .I1(n19646), .I2(n19645), .I3(n19644), .I4(n19643), .O(n19655)
         );
  AOI22S U22146 ( .A1(n20038), .A2(img[1923]), .B1(n19715), .B2(img[1795]), 
        .O(n19653) );
  AOI22S U22147 ( .A1(n19193), .A2(img[1667]), .B1(n13799), .B2(img[1539]), 
        .O(n19652) );
  AOI22S U22148 ( .A1(n13854), .A2(img[1411]), .B1(n19647), .B2(img[1283]), 
        .O(n19651) );
  AOI22S U22149 ( .A1(n13788), .A2(img[1155]), .B1(n13892), .B2(img[1027]), 
        .O(n19650) );
  AN4S U22150 ( .I1(n19653), .I2(n19652), .I3(n19651), .I4(n19650), .O(n19654)
         );
  ND2S U22151 ( .I1(n19655), .I2(n19654), .O(n19668) );
  AOI22S U22152 ( .A1(n19677), .A2(n20263), .B1(n13847), .B2(n19668), .O(
        n19659) );
  ND2S U22153 ( .I1(n19673), .I2(n21061), .O(n19658) );
  AOI22S U22154 ( .A1(n19666), .A2(n13804), .B1(n13846), .B2(n19701), .O(
        n19657) );
  AOI22S U22155 ( .A1(n19664), .A2(n13835), .B1(n13791), .B2(n19676), .O(
        n19656) );
  AN4S U22156 ( .I1(n19659), .I2(n19658), .I3(n19657), .I4(n19656), .O(n19694)
         );
  ND2S U22157 ( .I1(n19660), .I2(n19694), .O(n20320) );
  AOI22S U22158 ( .A1(n19663), .A2(n13839), .B1(n17875), .B2(n19662), .O(
        n19672) );
  AOI22S U22159 ( .A1(n19664), .A2(n19483), .B1(n20963), .B2(n19685), .O(
        n19671) );
  AOI22S U22160 ( .A1(n19666), .A2(n20124), .B1(n17762), .B2(n19665), .O(
        n19670) );
  AOI22S U22161 ( .A1(n19668), .A2(n13830), .B1(n17928), .B2(n19667), .O(
        n19669) );
  AN4S U22162 ( .I1(n19672), .I2(n19671), .I3(n19670), .I4(n19669), .O(n19683)
         );
  AOI22S U22163 ( .A1(n19673), .A2(n20439), .B1(n13847), .B2(n20315), .O(
        n19681) );
  ND2S U22164 ( .I1(n19674), .I2(n20580), .O(n19680) );
  AOI22S U22165 ( .A1(n19684), .A2(n13846), .B1(n13804), .B2(n19675), .O(
        n19679) );
  AOI22S U22166 ( .A1(n19677), .A2(n13791), .B1(n13793), .B2(n19676), .O(
        n19678) );
  AN4S U22167 ( .I1(n19681), .I2(n19680), .I3(n19679), .I4(n19678), .O(n19682)
         );
  ND2S U22168 ( .I1(n19683), .I2(n19682), .O(n19696) );
  AOI22S U22169 ( .A1(n20320), .A2(n20223), .B1(n20364), .B2(n19696), .O(
        n19699) );
  ND2S U22170 ( .I1(n19684), .I2(n13839), .O(n19687) );
  ND2S U22171 ( .I1(n19685), .I2(n17875), .O(n19686) );
  ND3S U22172 ( .I1(n19688), .I2(n19687), .I3(n19686), .O(n19692) );
  ND2S U22173 ( .I1(n19690), .I2(n19689), .O(n19691) );
  NR2 U22174 ( .I1(n19692), .I2(n19691), .O(n19693) );
  AO12 U22175 ( .B1(n19694), .B2(n19693), .A1(n19871), .O(n20321) );
  NR2 U22176 ( .I1(n13822), .I2(n20321), .O(n19695) );
  INV1S U22177 ( .I(n19695), .O(n19698) );
  ND2S U22178 ( .I1(n20062), .I2(n22932), .O(n19704) );
  ND2S U22179 ( .I1(n19701), .I2(n20366), .O(n19703) );
  AOI22S U22180 ( .A1(n20357), .A2(n20063), .B1(n19818), .B2(n19701), .O(
        n19702) );
  ND3 U22181 ( .I1(n19704), .I2(n19703), .I3(n19702), .O(n19705) );
  AOI22S U22182 ( .A1(n19745), .A2(n13839), .B1(n17875), .B2(n19744), .O(
        n19725) );
  AOI22S U22183 ( .A1(n19742), .A2(n21062), .B1(n20963), .B2(n19757), .O(
        n19724) );
  AOI22S U22184 ( .A1(n19743), .A2(n20613), .B1(n17762), .B2(n19755), .O(
        n19723) );
  AOI22S U22185 ( .A1(n13875), .A2(img[897]), .B1(n13797), .B2(img[769]), .O(
        n19714) );
  AOI22S U22186 ( .A1(n20102), .A2(img[641]), .B1(n19709), .B2(img[513]), .O(
        n19713) );
  AOI22S U22187 ( .A1(n19710), .A2(img[385]), .B1(n13836), .B2(img[257]), .O(
        n19712) );
  AOI22S U22188 ( .A1(n18819), .A2(img[129]), .B1(n20193), .B2(img[1]), .O(
        n19711) );
  AN4S U22189 ( .I1(n19714), .I2(n19713), .I3(n19712), .I4(n19711), .O(n19721)
         );
  AOI22S U22190 ( .A1(n13865), .A2(img[1921]), .B1(n19715), .B2(img[1793]), 
        .O(n19719) );
  AOI22S U22191 ( .A1(n17382), .A2(img[1665]), .B1(n13799), .B2(img[1537]), 
        .O(n19718) );
  AOI22S U22192 ( .A1(n13783), .A2(img[1409]), .B1(n15800), .B2(img[1281]), 
        .O(n19717) );
  AOI22S U22193 ( .A1(n18988), .A2(img[1153]), .B1(n13890), .B2(img[1025]), 
        .O(n19716) );
  AN4S U22194 ( .I1(n19719), .I2(n19718), .I3(n19717), .I4(n19716), .O(n19720)
         );
  ND2 U22195 ( .I1(n19721), .I2(n19720), .O(n19746) );
  AOI22S U22196 ( .A1(n19746), .A2(n13830), .B1(n17928), .B2(n19759), .O(
        n19722) );
  AN4S U22197 ( .I1(n19725), .I2(n19724), .I3(n19723), .I4(n19722), .O(n19731)
         );
  AOI22S U22198 ( .A1(n19756), .A2(n20439), .B1(n13847), .B2(n20324), .O(
        n19729) );
  ND2S U22199 ( .I1(n19758), .I2(n20150), .O(n19728) );
  AOI22S U22200 ( .A1(n19754), .A2(n13846), .B1(n13804), .B2(n19752), .O(
        n19727) );
  AOI22S U22201 ( .A1(n19747), .A2(n17938), .B1(n20406), .B2(n19753), .O(
        n19726) );
  AN4S U22202 ( .I1(n19729), .I2(n19728), .I3(n19727), .I4(n19726), .O(n19730)
         );
  ND2S U22203 ( .I1(n19731), .I2(n19730), .O(n19766) );
  AOI22S U22204 ( .A1(n19754), .A2(n13839), .B1(n17875), .B2(n19757), .O(
        n19735) );
  AOI22S U22205 ( .A1(n19759), .A2(n20963), .B1(n21062), .B2(n19745), .O(
        n19734) );
  AOI22S U22206 ( .A1(n19744), .A2(n20613), .B1(n17762), .B2(n19752), .O(
        n19733) );
  AOI22S U22207 ( .A1(n19755), .A2(n13830), .B1(n17928), .B2(n19758), .O(
        n19732) );
  AN4S U22208 ( .I1(n19735), .I2(n19734), .I3(n19733), .I4(n19732), .O(n19741)
         );
  AOI22S U22209 ( .A1(n19747), .A2(n20439), .B1(n13847), .B2(n19746), .O(
        n19739) );
  ND2S U22210 ( .I1(n19756), .I2(n21061), .O(n19738) );
  AOI22S U22211 ( .A1(n19743), .A2(n20620), .B1(n13846), .B2(n19770), .O(
        n19737) );
  AOI22S U22212 ( .A1(n19742), .A2(n19914), .B1(n13791), .B2(n19753), .O(
        n19736) );
  AOI22S U22213 ( .A1(n19766), .A2(n20364), .B1(n20223), .B2(n20329), .O(
        n19769) );
  AOI22S U22214 ( .A1(n19743), .A2(n20620), .B1(n13793), .B2(n19742), .O(
        n19751) );
  ND2S U22215 ( .I1(n19744), .I2(n20613), .O(n19750) );
  AOI22S U22216 ( .A1(n19746), .A2(n13847), .B1(n21062), .B2(n19745), .O(
        n19749) );
  AOI22S U22217 ( .A1(n19747), .A2(n20439), .B1(n13846), .B2(n19770), .O(
        n19748) );
  AN4S U22218 ( .I1(n19751), .I2(n19750), .I3(n19749), .I4(n19748), .O(n19765)
         );
  AOI22S U22219 ( .A1(n19753), .A2(n17938), .B1(n17762), .B2(n19752), .O(
        n19763) );
  AOI22S U22220 ( .A1(n19755), .A2(n13830), .B1(n13839), .B2(n19754), .O(
        n19762) );
  AOI22S U22221 ( .A1(n19757), .A2(n17875), .B1(n20629), .B2(n19756), .O(
        n19761) );
  AOI22S U22222 ( .A1(n19759), .A2(n20963), .B1(n17928), .B2(n19758), .O(
        n19760) );
  AN4S U22223 ( .I1(n19763), .I2(n19762), .I3(n19761), .I4(n19760), .O(n19764)
         );
  ND2S U22224 ( .I1(n19765), .I2(n19764), .O(n20330) );
  ND2S U22225 ( .I1(n20330), .I2(n20252), .O(n19768) );
  ND2 U22226 ( .I1(n19769), .I2(n13906), .O(n19775) );
  ND2S U22227 ( .I1(n20062), .I2(n13887), .O(n19773) );
  ND2S U22228 ( .I1(n19770), .I2(n20366), .O(n19772) );
  AOI22S U22229 ( .A1(n20343), .A2(n20063), .B1(n19818), .B2(n19770), .O(
        n19771) );
  ND3 U22230 ( .I1(n19773), .I2(n19772), .I3(n19771), .O(n19774) );
  OR2T U22231 ( .I1(n19775), .I2(n19774), .O(n23188) );
  AOI22S U22232 ( .A1(n20452), .A2(n20620), .B1(n20263), .B2(n20446), .O(
        n19779) );
  AOI22S U22233 ( .A1(n20454), .A2(n19914), .B1(n13847), .B2(n20453), .O(
        n19778) );
  AOI22S U22234 ( .A1(n20444), .A2(n13839), .B1(n13846), .B2(n20458), .O(
        n19777) );
  AOI22S U22235 ( .A1(n20457), .A2(n20187), .B1(n17938), .B2(n20442), .O(
        n19776) );
  AN4S U22236 ( .I1(n19779), .I2(n19778), .I3(n19777), .I4(n19776), .O(n19785)
         );
  AOI22S U22237 ( .A1(n20451), .A2(n20124), .B1(n17875), .B2(n20445), .O(
        n19783) );
  AOI22S U22238 ( .A1(n20456), .A2(n13830), .B1(n21062), .B2(n20443), .O(
        n19782) );
  AOI22S U22239 ( .A1(n20440), .A2(n20968), .B1(n17762), .B2(n20437), .O(
        n19781) );
  AOI22S U22240 ( .A1(n20455), .A2(n17928), .B1(n20969), .B2(n20441), .O(
        n19780) );
  AN4S U22241 ( .I1(n19783), .I2(n19782), .I3(n19781), .I4(n19780), .O(n19784)
         );
  ND2 U22242 ( .I1(n19785), .I2(n19784), .O(n19786) );
  MXL2HP U22243 ( .A(n23188), .B(n19786), .S(n13822), .OB(n21072) );
  INV2 U22244 ( .I(n21072), .O(n29462) );
  ND2S U22245 ( .I1(n29461), .I2(n29462), .O(n19850) );
  AOI22S U22246 ( .A1(n19835), .A2(n13839), .B1(n17875), .B2(n19827), .O(
        n19789) );
  AOI22S U22247 ( .A1(n19807), .A2(n20963), .B1(n19483), .B2(n19806), .O(
        n19830) );
  AOI22S U22248 ( .A1(n19824), .A2(n20613), .B1(n17762), .B2(n19840), .O(
        n19788) );
  AOI22S U22249 ( .A1(n19834), .A2(n13830), .B1(n17928), .B2(n19839), .O(
        n19787) );
  AN4S U22250 ( .I1(n19789), .I2(n19830), .I3(n19788), .I4(n19787), .O(n19805)
         );
  AOI22S U22251 ( .A1(n13875), .A2(img[896]), .B1(n13797), .B2(img[768]), .O(
        n19793) );
  AOI22S U22252 ( .A1(n19343), .A2(img[640]), .B1(n13859), .B2(img[512]), .O(
        n19792) );
  AOI22S U22253 ( .A1(n19949), .A2(img[384]), .B1(n17611), .B2(img[256]), .O(
        n19791) );
  AOI22S U22254 ( .A1(n17864), .A2(img[128]), .B1(n19950), .B2(img[0]), .O(
        n19790) );
  AN4S U22255 ( .I1(n19793), .I2(n19792), .I3(n19791), .I4(n19790), .O(n19799)
         );
  AOI22S U22256 ( .A1(n19215), .A2(img[1920]), .B1(n13794), .B2(img[1792]), 
        .O(n19797) );
  AOI22S U22257 ( .A1(n17382), .A2(img[1664]), .B1(n13798), .B2(img[1536]), 
        .O(n19796) );
  AOI22S U22258 ( .A1(n19856), .A2(img[1408]), .B1(n19955), .B2(img[1280]), 
        .O(n19795) );
  AOI22S U22259 ( .A1(n16037), .A2(img[1152]), .B1(n13890), .B2(img[1024]), 
        .O(n19794) );
  AN4S U22260 ( .I1(n19797), .I2(n19796), .I3(n19795), .I4(n19794), .O(n19798)
         );
  ND2S U22261 ( .I1(n19799), .I2(n19798), .O(n19836) );
  AOI22S U22262 ( .A1(n19825), .A2(n20439), .B1(n13847), .B2(n19836), .O(
        n19803) );
  ND2S U22263 ( .I1(n19833), .I2(n21061), .O(n19802) );
  AOI22S U22264 ( .A1(n19826), .A2(n13804), .B1(n13846), .B2(n19837), .O(
        n19801) );
  AOI22S U22265 ( .A1(n19828), .A2(n19914), .B1(n13791), .B2(n19838), .O(
        n19800) );
  AN4S U22266 ( .I1(n19803), .I2(n19802), .I3(n19801), .I4(n19800), .O(n19804)
         );
  ND2P U22267 ( .I1(n19805), .I2(n19804), .O(n20350) );
  AOI22S U22268 ( .A1(n19806), .A2(n13839), .B1(n17875), .B2(n19824), .O(
        n19811) );
  AOI22S U22269 ( .A1(n19828), .A2(n19483), .B1(n20963), .B2(n19827), .O(
        n19810) );
  AOI22S U22270 ( .A1(n19826), .A2(n20124), .B1(n17762), .B2(n19834), .O(
        n19809) );
  AOI22S U22271 ( .A1(n19836), .A2(n13830), .B1(n17928), .B2(n19807), .O(
        n19808) );
  AN4S U22272 ( .I1(n19811), .I2(n19810), .I3(n19809), .I4(n19808), .O(n19817)
         );
  AOI22S U22273 ( .A1(n19833), .A2(n20263), .B1(n13847), .B2(n20344), .O(
        n19815) );
  ND2S U22274 ( .I1(n19839), .I2(n20150), .O(n19814) );
  AOI22S U22275 ( .A1(n19835), .A2(n13846), .B1(n20438), .B2(n19840), .O(
        n19813) );
  AOI22S U22276 ( .A1(n19825), .A2(n17938), .B1(n13793), .B2(n19838), .O(
        n19812) );
  AN4S U22277 ( .I1(n19815), .I2(n19814), .I3(n19813), .I4(n19812), .O(n19816)
         );
  ND2S U22278 ( .I1(n19817), .I2(n19816), .O(n19823) );
  AOI22S U22279 ( .A1(n20350), .A2(n20223), .B1(n20364), .B2(n19823), .O(
        n19849) );
  ND2S U22280 ( .I1(n20062), .I2(n20345), .O(n19821) );
  ND2S U22281 ( .I1(n19837), .I2(n20366), .O(n19820) );
  AOI22S U22282 ( .A1(n20063), .A2(n20977), .B1(n19818), .B2(n19837), .O(
        n19819) );
  ND3 U22283 ( .I1(n19821), .I2(n19820), .I3(n19819), .O(n19822) );
  AOI12HS U22284 ( .B1(n19823), .B2(n20363), .A1(n19822), .O(n19848) );
  AOI22S U22285 ( .A1(n19825), .A2(n20263), .B1(n20613), .B2(n19824), .O(
        n19832) );
  ND2S U22286 ( .I1(n19826), .I2(n20620), .O(n19831) );
  AOI22S U22287 ( .A1(n19828), .A2(n19914), .B1(n17875), .B2(n19827), .O(
        n19829) );
  AN4S U22288 ( .I1(n19832), .I2(n19831), .I3(n19830), .I4(n19829), .O(n19846)
         );
  AOI22S U22289 ( .A1(n19834), .A2(n13830), .B1(n20629), .B2(n19833), .O(
        n19844) );
  AOI22S U22290 ( .A1(n19836), .A2(n13847), .B1(n13839), .B2(n19835), .O(
        n19843) );
  AOI22S U22291 ( .A1(n19838), .A2(n13791), .B1(n13846), .B2(n19837), .O(
        n19842) );
  AOI22S U22292 ( .A1(n19840), .A2(n17762), .B1(n17928), .B2(n19839), .O(
        n19841) );
  AN4S U22293 ( .I1(n19844), .I2(n19843), .I3(n19842), .I4(n19841), .O(n19845)
         );
  ND2S U22294 ( .I1(n19846), .I2(n19845), .O(n20351) );
  ND2S U22295 ( .I1(n20351), .I2(n20252), .O(n19847) );
  ND3P U22296 ( .I1(n19849), .I2(n19848), .I3(n19847), .O(n23187) );
  ND3S U22297 ( .I1(n19850), .I2(n23427), .I3(n21635), .O(n19913) );
  AOI22S U22298 ( .A1(n19326), .A2(img[898]), .B1(n13898), .B2(img[770]), .O(
        n19855) );
  AOI22S U22299 ( .A1(n13876), .A2(img[642]), .B1(n13859), .B2(img[514]), .O(
        n19854) );
  AOI22S U22300 ( .A1(n19949), .A2(img[386]), .B1(n17611), .B2(img[258]), .O(
        n19853) );
  AOI22S U22301 ( .A1(n20104), .A2(img[130]), .B1(n19950), .B2(img[2]), .O(
        n19852) );
  AN4S U22302 ( .I1(n19855), .I2(n19854), .I3(n19853), .I4(n19852), .O(n19862)
         );
  AOI22S U22303 ( .A1(n19215), .A2(img[1922]), .B1(n17561), .B2(img[1794]), 
        .O(n19860) );
  AOI22S U22304 ( .A1(n13823), .A2(img[1666]), .B1(n19182), .B2(img[1538]), 
        .O(n19859) );
  AOI22S U22305 ( .A1(n19856), .A2(img[1410]), .B1(n19955), .B2(img[1282]), 
        .O(n19858) );
  AOI22S U22306 ( .A1(n13788), .A2(img[1154]), .B1(n13890), .B2(img[1026]), 
        .O(n19857) );
  AN4S U22307 ( .I1(n19860), .I2(n19859), .I3(n19858), .I4(n19857), .O(n19861)
         );
  ND2S U22308 ( .I1(n19862), .I2(n19861), .O(n19886) );
  AOI22S U22309 ( .A1(n19895), .A2(n20263), .B1(n13847), .B2(n19886), .O(
        n19866) );
  ND2S U22310 ( .I1(n19891), .I2(n21061), .O(n19865) );
  AOI22S U22311 ( .A1(n19884), .A2(n20438), .B1(n13846), .B2(n19903), .O(
        n19864) );
  AOI22S U22312 ( .A1(n19881), .A2(n13835), .B1(n13791), .B2(n19896), .O(
        n19863) );
  AN4S U22313 ( .I1(n19866), .I2(n19865), .I3(n19864), .I4(n19863), .O(n19877)
         );
  AOI22S U22314 ( .A1(n19885), .A2(n20963), .B1(n19483), .B2(n19880), .O(
        n19875) );
  ND2S U22315 ( .I1(n19893), .I2(n13839), .O(n19868) );
  ND2S U22316 ( .I1(n19882), .I2(n17875), .O(n19867) );
  ND3S U22317 ( .I1(n19875), .I2(n19868), .I3(n19867), .O(n19870) );
  AOI22S U22318 ( .A1(n19879), .A2(n20613), .B1(n17762), .B2(n19894), .O(
        n19874) );
  AOI22S U22319 ( .A1(n19883), .A2(n13830), .B1(n17928), .B2(n19892), .O(
        n19873) );
  ND2S U22320 ( .I1(n19874), .I2(n19873), .O(n19869) );
  NR2 U22321 ( .I1(n19870), .I2(n19869), .O(n19872) );
  AO12 U22322 ( .B1(n19877), .B2(n19872), .A1(n19871), .O(n20340) );
  OR2 U22323 ( .I1(n13822), .I2(n20340), .O(n19911) );
  AOI22S U22324 ( .A1(n19893), .A2(n13839), .B1(n17875), .B2(n19882), .O(
        n19876) );
  AN4S U22325 ( .I1(n19876), .I2(n19875), .I3(n19874), .I4(n19873), .O(n19878)
         );
  ND2P U22326 ( .I1(n19878), .I2(n19877), .O(n20339) );
  AOI22S U22327 ( .A1(n19880), .A2(n13839), .B1(n17875), .B2(n19879), .O(
        n19890) );
  AOI22S U22328 ( .A1(n19882), .A2(n20963), .B1(n21062), .B2(n19881), .O(
        n19889) );
  AOI22S U22329 ( .A1(n19884), .A2(n20124), .B1(n17762), .B2(n19883), .O(
        n19888) );
  AOI22S U22330 ( .A1(n19886), .A2(n13830), .B1(n17928), .B2(n19885), .O(
        n19887) );
  AN4S U22331 ( .I1(n19890), .I2(n19889), .I3(n19888), .I4(n19887), .O(n19902)
         );
  AOI22S U22332 ( .A1(n20334), .A2(n13847), .B1(n20263), .B2(n19891), .O(
        n19900) );
  ND2S U22333 ( .I1(n19892), .I2(n20524), .O(n19899) );
  AOI22S U22334 ( .A1(n19894), .A2(n20620), .B1(n13846), .B2(n19893), .O(
        n19898) );
  AOI22S U22335 ( .A1(n19896), .A2(n19914), .B1(n13791), .B2(n19895), .O(
        n19897) );
  AN4S U22336 ( .I1(n19900), .I2(n19899), .I3(n19898), .I4(n19897), .O(n19901)
         );
  ND2S U22337 ( .I1(n19902), .I2(n19901), .O(n19908) );
  AOI22S U22338 ( .A1(n20339), .A2(n20223), .B1(n20364), .B2(n19908), .O(
        n19910) );
  ND2S U22339 ( .I1(n20062), .I2(n21225), .O(n19906) );
  ND2S U22340 ( .I1(n19903), .I2(n20366), .O(n19905) );
  ND3HT U22341 ( .I1(n19911), .I2(n19910), .I3(n19909), .O(n23186) );
  ND2S U22342 ( .I1(n20644), .I2(n23244), .O(n19912) );
  OAI112HS U22343 ( .C1(n23188), .C2(n29461), .A1(n19913), .B1(n19912), .O(
        n19927) );
  AOI22S U22344 ( .A1(n20477), .A2(n20620), .B1(n20439), .B2(n20476), .O(
        n19918) );
  AOI22S U22345 ( .A1(n20492), .A2(n19914), .B1(n13847), .B2(n20490), .O(
        n19917) );
  AOI22S U22346 ( .A1(n20475), .A2(n13839), .B1(n13846), .B2(n20484), .O(
        n19916) );
  AOI22S U22347 ( .A1(n20480), .A2(n20963), .B1(n13791), .B2(n20469), .O(
        n19915) );
  AN4S U22348 ( .I1(n19918), .I2(n19917), .I3(n19916), .I4(n19915), .O(n19924)
         );
  AOI22S U22349 ( .A1(n20489), .A2(n20613), .B1(n17875), .B2(n20474), .O(
        n19922) );
  AOI22S U22350 ( .A1(n20485), .A2(n13830), .B1(n21062), .B2(n20471), .O(
        n19921) );
  AOI22S U22351 ( .A1(n20468), .A2(n18040), .B1(n17762), .B2(n20481), .O(
        n19920) );
  AOI22S U22352 ( .A1(n20491), .A2(n17928), .B1(n20969), .B2(n20470), .O(
        n19919) );
  AN4S U22353 ( .I1(n19922), .I2(n19921), .I3(n19920), .I4(n19919), .O(n19923)
         );
  MXL2HP U22354 ( .A(n23186), .B(n19925), .S(n13822), .OB(n21076) );
  ND2S U22355 ( .I1(n29484), .I2(n29483), .O(n19926) );
  OAI112HS U22356 ( .C1(n20503), .C2(n21079), .A1(n19927), .B1(n19926), .O(
        n20183) );
  INV1S U22357 ( .I(n20942), .O(n19928) );
  ND2S U22358 ( .I1(n19928), .I2(n21811), .O(n20182) );
  INV1S U22359 ( .I(n19929), .O(n20574) );
  MOAI1S U22360 ( .A1(n13947), .A2(n20574), .B1(n20569), .B2(n14174), .O(
        n19933) );
  INV1S U22361 ( .I(n19930), .O(n20586) );
  MOAI1S U22362 ( .A1(n13927), .A2(n20586), .B1(n20577), .B2(n19931), .O(
        n19932) );
  NR2 U22363 ( .I1(n19933), .I2(n19932), .O(n19936) );
  AOI22S U22364 ( .A1(n20595), .A2(n20439), .B1(n13835), .B2(n20581), .O(
        n19935) );
  AOI22S U22365 ( .A1(n20578), .A2(n13847), .B1(n13839), .B2(n20593), .O(
        n19934) );
  ND2S U22366 ( .I1(n20579), .I2(n17928), .O(n19938) );
  ND2S U22367 ( .I1(n20594), .I2(n20620), .O(n19937) );
  ND3S U22368 ( .I1(n19938), .I2(n19937), .I3(n13822), .O(n19941) );
  INV1S U22369 ( .I(n19939), .O(n20589) );
  MOAI1S U22370 ( .A1(n13844), .A2(n20589), .B1(n20570), .B2(n17762), .O(
        n19940) );
  NR2 U22371 ( .I1(n19941), .I2(n19940), .O(n19944) );
  AOI22S U22372 ( .A1(n20592), .A2(n17875), .B1(n13830), .B2(n20573), .O(
        n19943) );
  AOI22S U22373 ( .A1(n20588), .A2(n19483), .B1(n20629), .B2(n20585), .O(
        n19942) );
  ND3S U22374 ( .I1(n19944), .I2(n19943), .I3(n19942), .O(n20011) );
  AOI22S U22375 ( .A1(n19983), .A2(n13839), .B1(n17875), .B2(n20000), .O(
        n19948) );
  AOI22S U22376 ( .A1(n19997), .A2(n20963), .B1(n21062), .B2(n19994), .O(
        n19947) );
  AOI22S U22377 ( .A1(n19999), .A2(n20613), .B1(n17762), .B2(n19985), .O(
        n19946) );
  AOI22S U22378 ( .A1(n20001), .A2(n13830), .B1(n17928), .B2(n19995), .O(
        n19945) );
  AN4S U22379 ( .I1(n19948), .I2(n19947), .I3(n19946), .I4(n19945), .O(n19968)
         );
  AOI22S U22380 ( .A1(n13875), .A2(img[902]), .B1(n13837), .B2(img[774]), .O(
        n19954) );
  AOI22S U22381 ( .A1(n13785), .A2(img[646]), .B1(n13879), .B2(img[518]), .O(
        n19953) );
  AOI22S U22382 ( .A1(n19949), .A2(img[390]), .B1(n17611), .B2(img[262]), .O(
        n19952) );
  AOI22S U22383 ( .A1(n17778), .A2(img[134]), .B1(n19950), .B2(img[6]), .O(
        n19951) );
  AN4S U22384 ( .I1(n19954), .I2(n19953), .I3(n19952), .I4(n19951), .O(n19962)
         );
  AOI22S U22385 ( .A1(n15809), .A2(img[1926]), .B1(n19416), .B2(img[1798]), 
        .O(n19960) );
  AOI22S U22386 ( .A1(n15630), .A2(img[1670]), .B1(n19182), .B2(img[1542]), 
        .O(n19959) );
  AOI22S U22387 ( .A1(n18778), .A2(img[1414]), .B1(n19955), .B2(img[1286]), 
        .O(n19958) );
  AOI22S U22388 ( .A1(n19649), .A2(img[1158]), .B1(n13880), .B2(img[1030]), 
        .O(n19957) );
  AN4S U22389 ( .I1(n19960), .I2(n19959), .I3(n19958), .I4(n19957), .O(n19961)
         );
  ND2S U22390 ( .I1(n19962), .I2(n19961), .O(n19984) );
  AOI22S U22391 ( .A1(n19998), .A2(n20439), .B1(n13847), .B2(n19984), .O(
        n19966) );
  ND2S U22392 ( .I1(n19996), .I2(n20150), .O(n19965) );
  AOI22S U22393 ( .A1(n19989), .A2(n13804), .B1(n13846), .B2(n19987), .O(
        n19964) );
  AOI22S U22394 ( .A1(n19986), .A2(n19914), .B1(n13791), .B2(n19988), .O(
        n19963) );
  AN4S U22395 ( .I1(n19966), .I2(n19965), .I3(n19964), .I4(n19963), .O(n19967)
         );
  AOI22S U22396 ( .A1(n19994), .A2(n13839), .B1(n17875), .B2(n19999), .O(
        n19972) );
  AOI22S U22397 ( .A1(n19986), .A2(n21062), .B1(n20963), .B2(n20000), .O(
        n19971) );
  AOI22S U22398 ( .A1(n19989), .A2(n20613), .B1(n17762), .B2(n20001), .O(
        n19970) );
  AOI22S U22399 ( .A1(n19984), .A2(n13830), .B1(n17928), .B2(n19997), .O(
        n19969) );
  AN4S U22400 ( .I1(n19972), .I2(n19971), .I3(n19970), .I4(n19969), .O(n19978)
         );
  AOI22S U22401 ( .A1(n19996), .A2(n20439), .B1(n13847), .B2(n20293), .O(
        n19976) );
  ND2S U22402 ( .I1(n19995), .I2(n20524), .O(n19975) );
  AOI22S U22403 ( .A1(n19983), .A2(n13846), .B1(n20438), .B2(n19985), .O(
        n19974) );
  AOI22S U22404 ( .A1(n19998), .A2(n13791), .B1(n13793), .B2(n19988), .O(
        n19973) );
  AN4S U22405 ( .I1(n19976), .I2(n19975), .I3(n19974), .I4(n19973), .O(n19977)
         );
  ND2S U22406 ( .I1(n19978), .I2(n19977), .O(n19979) );
  AOI22S U22407 ( .A1(n20298), .A2(n20223), .B1(n20364), .B2(n19979), .O(
        n20010) );
  ND2S U22408 ( .I1(n20062), .I2(n21254), .O(n19980) );
  AOI22S U22409 ( .A1(n19984), .A2(n13847), .B1(n13839), .B2(n19983), .O(
        n19993) );
  ND2S U22410 ( .I1(n19985), .I2(n17762), .O(n19992) );
  AOI22S U22411 ( .A1(n19987), .A2(n13846), .B1(n13793), .B2(n19986), .O(
        n19991) );
  AOI22S U22412 ( .A1(n19989), .A2(n13804), .B1(n17938), .B2(n19988), .O(
        n19990) );
  AN4S U22413 ( .I1(n19993), .I2(n19992), .I3(n19991), .I4(n19990), .O(n20007)
         );
  AOI22S U22414 ( .A1(n19995), .A2(n17928), .B1(n21062), .B2(n19994), .O(
        n20005) );
  AOI22S U22415 ( .A1(n19997), .A2(n20963), .B1(n20560), .B2(n19996), .O(
        n20004) );
  AOI22S U22416 ( .A1(n19999), .A2(n20613), .B1(n20439), .B2(n19998), .O(
        n20003) );
  AOI22S U22417 ( .A1(n20001), .A2(n13830), .B1(n17875), .B2(n20000), .O(
        n20002) );
  AN4S U22418 ( .I1(n20005), .I2(n20004), .I3(n20003), .I4(n20002), .O(n20006)
         );
  ND2S U22419 ( .I1(n20007), .I2(n20006), .O(n20299) );
  ND2S U22420 ( .I1(n20299), .I2(n20252), .O(n20008) );
  ND3P U22421 ( .I1(n20010), .I2(n20009), .I3(n20008), .O(n23179) );
  OR2P U22422 ( .I1(n13822), .I2(n23179), .O(n20949) );
  OAI12HP U22423 ( .B1(n20012), .B2(n20011), .A1(n20949), .O(n21088) );
  ND2S U22424 ( .I1(n29505), .I2(n29503), .O(n20186) );
  INV1S U22425 ( .I(n20013), .O(n20556) );
  MOAI1S U22426 ( .A1(n13947), .A2(n20556), .B1(n20551), .B2(n20963), .O(
        n20016) );
  INV1S U22427 ( .I(n20540), .O(n20014) );
  MOAI1S U22428 ( .A1(n13927), .A2(n20014), .B1(n20557), .B2(n20613), .O(
        n20015) );
  NR2 U22429 ( .I1(n20016), .I2(n20015), .O(n20019) );
  AOI22S U22430 ( .A1(n20546), .A2(n20439), .B1(n13793), .B2(n20561), .O(
        n20018) );
  AOI22S U22431 ( .A1(n20558), .A2(n13847), .B1(n13839), .B2(n20544), .O(
        n20017) );
  ND3S U22432 ( .I1(n20019), .I2(n20018), .I3(n20017), .O(n20098) );
  ND2S U22433 ( .I1(n20559), .I2(n17928), .O(n20021) );
  ND2S U22434 ( .I1(n20545), .I2(n13804), .O(n20020) );
  ND3S U22435 ( .I1(n20021), .I2(n20020), .I3(n13822), .O(n20024) );
  INV1S U22436 ( .I(n20541), .O(n20022) );
  MOAI1S U22437 ( .A1(n13844), .A2(n20022), .B1(n20552), .B2(n17762), .O(
        n20023) );
  NR2 U22438 ( .I1(n20024), .I2(n20023), .O(n20027) );
  AOI22S U22439 ( .A1(n20543), .A2(n17875), .B1(n13830), .B2(n20555), .O(
        n20026) );
  AOI22S U22440 ( .A1(n20542), .A2(n19483), .B1(n20629), .B2(n20539), .O(
        n20025) );
  ND3 U22441 ( .I1(n20027), .I2(n20026), .I3(n20025), .O(n20097) );
  AOI22S U22442 ( .A1(n20072), .A2(n13839), .B1(n17875), .B2(n20084), .O(
        n20031) );
  AOI22S U22443 ( .A1(n20069), .A2(n20963), .B1(n21062), .B2(n20074), .O(
        n20030) );
  AOI22S U22444 ( .A1(n20087), .A2(n20613), .B1(n17762), .B2(n20075), .O(
        n20029) );
  AOI22S U22445 ( .A1(n20085), .A2(n13830), .B1(n17928), .B2(n20082), .O(
        n20028) );
  AN4S U22446 ( .I1(n20031), .I2(n20030), .I3(n20029), .I4(n20028), .O(n20051)
         );
  AOI22S U22447 ( .A1(n17835), .A2(img[901]), .B1(n13898), .B2(img[773]), .O(
        n20037) );
  AOI22S U22448 ( .A1(n20032), .A2(img[645]), .B1(n13858), .B2(img[517]), .O(
        n20036) );
  AOI22S U22449 ( .A1(n13800), .A2(img[389]), .B1(n19388), .B2(img[261]), .O(
        n20035) );
  AOI22S U22450 ( .A1(n18958), .A2(img[133]), .B1(n20033), .B2(img[5]), .O(
        n20034) );
  AN4S U22451 ( .I1(n20037), .I2(n20036), .I3(n20035), .I4(n20034), .O(n20045)
         );
  AOI22S U22452 ( .A1(n20038), .A2(img[1925]), .B1(n13796), .B2(img[1797]), 
        .O(n20043) );
  AOI22S U22453 ( .A1(n18837), .A2(img[1669]), .B1(n13799), .B2(img[1541]), 
        .O(n20042) );
  AOI22S U22454 ( .A1(n17359), .A2(img[1413]), .B1(n20039), .B2(img[1285]), 
        .O(n20041) );
  AOI22S U22455 ( .A1(n13788), .A2(img[1157]), .B1(n13880), .B2(img[1029]), 
        .O(n20040) );
  AN4S U22456 ( .I1(n20043), .I2(n20042), .I3(n20041), .I4(n20040), .O(n20044)
         );
  ND2S U22457 ( .I1(n20045), .I2(n20044), .O(n20071) );
  AOI22S U22458 ( .A1(n20083), .A2(n20263), .B1(n13847), .B2(n20071), .O(
        n20049) );
  ND2S U22459 ( .I1(n20081), .I2(n21061), .O(n20048) );
  AOI22S U22460 ( .A1(n20070), .A2(n13804), .B1(n13846), .B2(n20080), .O(
        n20047) );
  AOI22S U22461 ( .A1(n20086), .A2(n19914), .B1(n13791), .B2(n20073), .O(
        n20046) );
  AN4S U22462 ( .I1(n20049), .I2(n20048), .I3(n20047), .I4(n20046), .O(n20050)
         );
  ND2 U22463 ( .I1(n20051), .I2(n20050), .O(n20308) );
  AOI22S U22464 ( .A1(n20074), .A2(n13839), .B1(n17875), .B2(n20087), .O(
        n20055) );
  AOI22S U22465 ( .A1(n20086), .A2(n19483), .B1(n20963), .B2(n20084), .O(
        n20054) );
  AOI22S U22466 ( .A1(n20070), .A2(n20613), .B1(n17762), .B2(n20085), .O(
        n20053) );
  AOI22S U22467 ( .A1(n20071), .A2(n13830), .B1(n17928), .B2(n20069), .O(
        n20052) );
  AN4S U22468 ( .I1(n20055), .I2(n20054), .I3(n20053), .I4(n20052), .O(n20061)
         );
  AOI22S U22469 ( .A1(n20081), .A2(n20439), .B1(n13847), .B2(n20303), .O(
        n20059) );
  ND2S U22470 ( .I1(n20082), .I2(n20150), .O(n20058) );
  AOI22S U22471 ( .A1(n20072), .A2(n13846), .B1(n20438), .B2(n20075), .O(
        n20057) );
  AOI22S U22472 ( .A1(n20083), .A2(n13791), .B1(n13793), .B2(n20073), .O(
        n20056) );
  AN4S U22473 ( .I1(n20059), .I2(n20058), .I3(n20057), .I4(n20056), .O(n20060)
         );
  ND2S U22474 ( .I1(n20061), .I2(n20060), .O(n20068) );
  AOI22S U22475 ( .A1(n20308), .A2(n20223), .B1(n20364), .B2(n20068), .O(
        n20096) );
  ND2S U22476 ( .I1(n20062), .I2(n21245), .O(n20066) );
  ND2S U22477 ( .I1(n20080), .I2(n20366), .O(n20065) );
  AOI22S U22478 ( .A1(n20688), .A2(n20063), .B1(n19818), .B2(n20080), .O(
        n20064) );
  ND3S U22479 ( .I1(n20066), .I2(n20065), .I3(n20064), .O(n20067) );
  AOI12HS U22480 ( .B1(n20068), .B2(n20363), .A1(n20067), .O(n20095) );
  AOI22S U22481 ( .A1(n20070), .A2(n13804), .B1(n20963), .B2(n20069), .O(
        n20079) );
  ND2S U22482 ( .I1(n20071), .I2(n13847), .O(n20078) );
  AOI22S U22483 ( .A1(n20073), .A2(n13791), .B1(n13839), .B2(n20072), .O(
        n20077) );
  AOI22S U22484 ( .A1(n20075), .A2(n17762), .B1(n19483), .B2(n20074), .O(
        n20076) );
  AN4S U22485 ( .I1(n20079), .I2(n20078), .I3(n20077), .I4(n20076), .O(n20093)
         );
  AOI22S U22486 ( .A1(n20081), .A2(n20968), .B1(n13846), .B2(n20080), .O(
        n20091) );
  AOI22S U22487 ( .A1(n20083), .A2(n20263), .B1(n17928), .B2(n20082), .O(
        n20090) );
  AOI22S U22488 ( .A1(n20085), .A2(n13830), .B1(n17875), .B2(n20084), .O(
        n20089) );
  AOI22S U22489 ( .A1(n20087), .A2(n20613), .B1(n13793), .B2(n20086), .O(
        n20088) );
  AN4S U22490 ( .I1(n20091), .I2(n20090), .I3(n20089), .I4(n20088), .O(n20092)
         );
  ND2S U22491 ( .I1(n20093), .I2(n20092), .O(n20309) );
  ND2S U22492 ( .I1(n20309), .I2(n20252), .O(n20094) );
  OAI12HP U22493 ( .B1(n20098), .B2(n20097), .A1(n21000), .O(n21081) );
  ND2S U22494 ( .I1(n26015), .I2(n21595), .O(n20185) );
  AOI22S U22495 ( .A1(n20129), .A2(n13839), .B1(n17875), .B2(n20123), .O(
        n20147) );
  ND2S U22496 ( .I1(n20140), .I2(n17762), .O(n20101) );
  AOI22S U22497 ( .A1(n20139), .A2(n20187), .B1(n20406), .B2(n20154), .O(
        n20100) );
  AOI22S U22498 ( .A1(n20152), .A2(n20620), .B1(n13791), .B2(n20153), .O(
        n20099) );
  AN4S U22499 ( .I1(n20147), .I2(n20101), .I3(n20100), .I4(n20099), .O(n20122)
         );
  AOI22S U22500 ( .A1(n20141), .A2(n20124), .B1(n13846), .B2(n20163), .O(
        n20120) );
  AOI22S U22501 ( .A1(n20143), .A2(n13830), .B1(n20439), .B2(n20149), .O(
        n20119) );
  AOI22S U22502 ( .A1(n20151), .A2(n18040), .B1(n19483), .B2(n20138), .O(
        n20118) );
  AOI22S U22503 ( .A1(n13875), .A2(img[900]), .B1(n13797), .B2(img[772]), .O(
        n20108) );
  AOI22S U22504 ( .A1(n20102), .A2(img[644]), .B1(n13858), .B2(img[516]), .O(
        n20107) );
  AOI22S U22505 ( .A1(n19710), .A2(img[388]), .B1(n20103), .B2(img[260]), .O(
        n20106) );
  AOI22S U22506 ( .A1(n17335), .A2(img[132]), .B1(n20193), .B2(img[4]), .O(
        n20105) );
  AN4S U22507 ( .I1(n20108), .I2(n20107), .I3(n20106), .I4(n20105), .O(n20116)
         );
  AOI22S U22508 ( .A1(n19036), .A2(img[1924]), .B1(n19416), .B2(img[1796]), 
        .O(n20114) );
  AOI22S U22509 ( .A1(n20109), .A2(img[1668]), .B1(n13845), .B2(img[1540]), 
        .O(n20113) );
  AOI22S U22510 ( .A1(n13783), .A2(img[1412]), .B1(n15800), .B2(img[1284]), 
        .O(n20112) );
  AOI22S U22511 ( .A1(n16515), .A2(img[1156]), .B1(n16048), .B2(img[1028]), 
        .O(n20111) );
  AN4S U22512 ( .I1(n20114), .I2(n20113), .I3(n20112), .I4(n20111), .O(n20115)
         );
  ND2 U22513 ( .I1(n20116), .I2(n20115), .O(n20148) );
  AOI22S U22514 ( .A1(n20148), .A2(n13847), .B1(n17928), .B2(n20142), .O(
        n20117) );
  AN4S U22515 ( .I1(n20120), .I2(n20119), .I3(n20118), .I4(n20117), .O(n20121)
         );
  ND2S U22516 ( .I1(n20122), .I2(n20121), .O(n20374) );
  ND2S U22517 ( .I1(n20374), .I2(n20252), .O(n20137) );
  AOI22S U22518 ( .A1(n20138), .A2(n13839), .B1(n17875), .B2(n20141), .O(
        n20128) );
  AOI22S U22519 ( .A1(n20154), .A2(n21062), .B1(n20963), .B2(n20123), .O(
        n20127) );
  AOI22S U22520 ( .A1(n20152), .A2(n20124), .B1(n17762), .B2(n20143), .O(
        n20126) );
  AOI22S U22521 ( .A1(n20148), .A2(n13830), .B1(n17928), .B2(n20139), .O(
        n20125) );
  AN4S U22522 ( .I1(n20128), .I2(n20127), .I3(n20126), .I4(n20125), .O(n20135)
         );
  AOI22S U22523 ( .A1(n20151), .A2(n20439), .B1(n13847), .B2(n20365), .O(
        n20133) );
  ND2S U22524 ( .I1(n20142), .I2(n20560), .O(n20132) );
  AOI22S U22525 ( .A1(n20129), .A2(n13846), .B1(n20438), .B2(n20140), .O(
        n20131) );
  AOI22S U22526 ( .A1(n20149), .A2(n17938), .B1(n13793), .B2(n20153), .O(
        n20130) );
  AN4S U22527 ( .I1(n20133), .I2(n20132), .I3(n20131), .I4(n20130), .O(n20134)
         );
  ND2S U22528 ( .I1(n20135), .I2(n20134), .O(n20161) );
  AOI22S U22529 ( .A1(n20139), .A2(n20963), .B1(n21062), .B2(n20138), .O(
        n20146) );
  AOI22S U22530 ( .A1(n20141), .A2(n20613), .B1(n17762), .B2(n20140), .O(
        n20145) );
  AOI22S U22531 ( .A1(n20143), .A2(n13830), .B1(n17928), .B2(n20142), .O(
        n20144) );
  AN4S U22532 ( .I1(n20147), .I2(n20146), .I3(n20145), .I4(n20144), .O(n20160)
         );
  AOI22S U22533 ( .A1(n20149), .A2(n20439), .B1(n13847), .B2(n20148), .O(
        n20158) );
  ND2S U22534 ( .I1(n20151), .I2(n20150), .O(n20157) );
  AOI22S U22535 ( .A1(n20152), .A2(n13804), .B1(n13846), .B2(n20163), .O(
        n20156) );
  AOI22S U22536 ( .A1(n20154), .A2(n19914), .B1(n13791), .B2(n20153), .O(
        n20155) );
  AN4S U22537 ( .I1(n20158), .I2(n20157), .I3(n20156), .I4(n20155), .O(n20159)
         );
  AOI22S U22538 ( .A1(n20372), .A2(n20223), .B1(n20364), .B2(n20161), .O(
        n20162) );
  ND2 U22539 ( .I1(n13936), .I2(n20162), .O(n20168) );
  ND2S U22540 ( .I1(n20163), .I2(n20366), .O(n20166) );
  ND2S U22541 ( .I1(n20740), .I2(n18142), .O(n20165) );
  ND2S U22542 ( .I1(n20163), .I2(n19818), .O(n20164) );
  ND3 U22543 ( .I1(n20166), .I2(n20165), .I3(n20164), .O(n20167) );
  AOI22S U22544 ( .A1(n20520), .A2(n20620), .B1(n20263), .B2(n20514), .O(
        n20172) );
  AOI22S U22545 ( .A1(n20522), .A2(n13793), .B1(n13847), .B2(n20521), .O(
        n20171) );
  AOI22S U22546 ( .A1(n20512), .A2(n13839), .B1(n13846), .B2(n20527), .O(
        n20170) );
  AOI22S U22547 ( .A1(n20526), .A2(n20963), .B1(n13791), .B2(n20510), .O(
        n20169) );
  AN4S U22548 ( .I1(n20172), .I2(n20171), .I3(n20170), .I4(n20169), .O(n20178)
         );
  AOI22S U22549 ( .A1(n20519), .A2(n20124), .B1(n17875), .B2(n20513), .O(
        n20176) );
  AOI22S U22550 ( .A1(n20525), .A2(n13830), .B1(n19483), .B2(n20511), .O(
        n20175) );
  AOI22S U22551 ( .A1(n20508), .A2(n20560), .B1(n17762), .B2(n20507), .O(
        n20174) );
  AOI22S U22552 ( .A1(n20523), .A2(n17928), .B1(n20969), .B2(n20509), .O(
        n20173) );
  AN4S U22553 ( .I1(n20176), .I2(n20175), .I3(n20174), .I4(n20173), .O(n20177)
         );
  ND2 U22554 ( .I1(n20178), .I2(n20177), .O(n20179) );
  MXL2HP U22555 ( .A(n23184), .B(n20179), .S(n13822), .OB(n21023) );
  INV2 U22556 ( .I(n21023), .O(n28533) );
  ND2S U22557 ( .I1(n21611), .I2(n28533), .O(n20180) );
  ND3 U22558 ( .I1(n20186), .I2(n20185), .I3(n20180), .O(n20181) );
  AOI12HS U22559 ( .B1(n20183), .B2(n20182), .A1(n20181), .O(n20279) );
  OAI22S U22560 ( .A1(n23184), .A2(n21611), .B1(n13814), .B2(n21000), .O(
        n20184) );
  ND3S U22561 ( .I1(n20186), .I2(n20185), .I3(n20184), .O(n20258) );
  INV1S U22562 ( .I(n20949), .O(n21006) );
  ND2S U22563 ( .I1(n21006), .I2(n21804), .O(n20257) );
  AOI22S U22564 ( .A1(n20233), .A2(n13839), .B1(n17875), .B2(n20234), .O(
        n20190) );
  AOI22S U22565 ( .A1(n20212), .A2(n20187), .B1(n19483), .B2(n20211), .O(
        n20248) );
  AOI22S U22566 ( .A1(n20241), .A2(n20613), .B1(n17762), .B2(n20229), .O(
        n20189) );
  AOI22S U22567 ( .A1(n20243), .A2(n13830), .B1(n17928), .B2(n20245), .O(
        n20188) );
  AOI22S U22568 ( .A1(n19252), .A2(img[903]), .B1(n13898), .B2(img[775]), .O(
        n20197) );
  AOI22S U22569 ( .A1(n13876), .A2(img[647]), .B1(n13858), .B2(img[519]), .O(
        n20196) );
  AOI22S U22570 ( .A1(n20192), .A2(img[391]), .B1(n13836), .B2(img[263]), .O(
        n20195) );
  AOI22S U22571 ( .A1(n17886), .A2(img[135]), .B1(n20193), .B2(img[7]), .O(
        n20194) );
  AN4S U22572 ( .I1(n20197), .I2(n20196), .I3(n20195), .I4(n20194), .O(n20204)
         );
  AOI22S U22573 ( .A1(n19036), .A2(img[1927]), .B1(n18201), .B2(img[1799]), 
        .O(n20202) );
  AOI22S U22574 ( .A1(n13823), .A2(img[1671]), .B1(n18751), .B2(img[1543]), 
        .O(n20201) );
  AOI22S U22575 ( .A1(n18778), .A2(img[1415]), .B1(n20198), .B2(img[1287]), 
        .O(n20200) );
  AOI22S U22576 ( .A1(n18946), .A2(img[1159]), .B1(n15653), .B2(img[1031]), 
        .O(n20199) );
  AN4S U22577 ( .I1(n20202), .I2(n20201), .I3(n20200), .I4(n20199), .O(n20203)
         );
  ND2S U22578 ( .I1(n20204), .I2(n20203), .O(n20230) );
  AOI22S U22579 ( .A1(n20235), .A2(n20263), .B1(n13847), .B2(n20230), .O(
        n20208) );
  ND2S U22580 ( .I1(n20242), .I2(n20580), .O(n20207) );
  AOI22S U22581 ( .A1(n20231), .A2(n20620), .B1(n13846), .B2(n20244), .O(
        n20206) );
  AOI22S U22582 ( .A1(n20240), .A2(n13793), .B1(n13791), .B2(n20232), .O(
        n20205) );
  AN4S U22583 ( .I1(n20208), .I2(n20207), .I3(n20206), .I4(n20205), .O(n20209)
         );
  ND2 U22584 ( .I1(n20210), .I2(n20209), .O(n20286) );
  AOI22S U22585 ( .A1(n20211), .A2(n13839), .B1(n17875), .B2(n20241), .O(
        n20216) );
  AOI22S U22586 ( .A1(n20240), .A2(n19483), .B1(n20187), .B2(n20234), .O(
        n20215) );
  AOI22S U22587 ( .A1(n20231), .A2(n20124), .B1(n17762), .B2(n20243), .O(
        n20214) );
  AOI22S U22588 ( .A1(n20230), .A2(n13830), .B1(n17928), .B2(n20212), .O(
        n20213) );
  AN4S U22589 ( .I1(n20216), .I2(n20215), .I3(n20214), .I4(n20213), .O(n20222)
         );
  AOI22S U22590 ( .A1(n20242), .A2(n20439), .B1(n13847), .B2(n20281), .O(
        n20220) );
  ND2S U22591 ( .I1(n20245), .I2(n21061), .O(n20219) );
  AOI22S U22592 ( .A1(n20233), .A2(n13846), .B1(n20438), .B2(n20229), .O(
        n20218) );
  AOI22S U22593 ( .A1(n20235), .A2(n13791), .B1(n20406), .B2(n20232), .O(
        n20217) );
  AN4S U22594 ( .I1(n20220), .I2(n20219), .I3(n20218), .I4(n20217), .O(n20221)
         );
  AOI22S U22595 ( .A1(n20286), .A2(n20223), .B1(n16188), .B2(n20228), .O(
        n20255) );
  ND2 U22596 ( .I1(n21669), .I2(n18142), .O(n20225) );
  AOI12HS U22597 ( .B1(n20228), .B2(n20363), .A1(n20227), .O(n20254) );
  AOI22S U22598 ( .A1(n20230), .A2(n13847), .B1(n17762), .B2(n20229), .O(
        n20239) );
  ND2S U22599 ( .I1(n20231), .I2(n20620), .O(n20238) );
  AOI22S U22600 ( .A1(n20233), .A2(n13839), .B1(n13791), .B2(n20232), .O(
        n20237) );
  AOI22S U22601 ( .A1(n20235), .A2(n20263), .B1(n17875), .B2(n20234), .O(
        n20236) );
  AN4S U22602 ( .I1(n20239), .I2(n20238), .I3(n20237), .I4(n20236), .O(n20251)
         );
  AOI22S U22603 ( .A1(n20241), .A2(n20613), .B1(n13793), .B2(n20240), .O(
        n20249) );
  AOI22S U22604 ( .A1(n20243), .A2(n13830), .B1(n18040), .B2(n20242), .O(
        n20247) );
  AOI22S U22605 ( .A1(n20245), .A2(n17928), .B1(n13846), .B2(n20244), .O(
        n20246) );
  AN4S U22606 ( .I1(n20249), .I2(n20248), .I3(n20247), .I4(n20246), .O(n20250)
         );
  ND2S U22607 ( .I1(n20251), .I2(n20250), .O(n20287) );
  ND3P U22608 ( .I1(n20255), .I2(n20254), .I3(n20253), .O(n23178) );
  OR2 U22609 ( .I1(n23178), .I2(n21467), .O(n20256) );
  ND3S U22610 ( .I1(n20258), .I2(n20257), .I3(n20256), .O(n20278) );
  INV1S U22611 ( .I(n20259), .O(n20625) );
  MOAI1S U22612 ( .A1(n13947), .A2(n20625), .B1(n20619), .B2(n14174), .O(
        n20262) );
  INV1S U22613 ( .I(n20607), .O(n20260) );
  MOAI1S U22614 ( .A1(n13927), .A2(n20260), .B1(n20626), .B2(n20613), .O(
        n20261) );
  NR2 U22615 ( .I1(n20262), .I2(n20261), .O(n20266) );
  AOI22S U22616 ( .A1(n20614), .A2(n20263), .B1(n20406), .B2(n20630), .O(
        n20265) );
  AOI22S U22617 ( .A1(n20627), .A2(n13847), .B1(n13839), .B2(n20611), .O(
        n20264) );
  ND2S U22618 ( .I1(n20628), .I2(n17928), .O(n20268) );
  ND2S U22619 ( .I1(n20612), .I2(n20620), .O(n20267) );
  ND3S U22620 ( .I1(n20268), .I2(n20267), .I3(n13822), .O(n20271) );
  INV1S U22621 ( .I(n20608), .O(n20269) );
  MOAI1S U22622 ( .A1(n13844), .A2(n20269), .B1(n20621), .B2(n17762), .O(
        n20270) );
  NR2 U22623 ( .I1(n20271), .I2(n20270), .O(n20274) );
  AOI22S U22624 ( .A1(n20610), .A2(n17875), .B1(n13830), .B2(n20624), .O(
        n20273) );
  AOI22S U22625 ( .A1(n20609), .A2(n19483), .B1(n20629), .B2(n20606), .O(
        n20272) );
  OR2T U22626 ( .I1(n13822), .I2(n23178), .O(n20948) );
  OAI12HP U22627 ( .B1(n20276), .B2(n20275), .A1(n20948), .O(n21085) );
  ND2S U22628 ( .I1(n23848), .I2(n21467), .O(n20277) );
  OA12P U22629 ( .B1(n20279), .B2(n20278), .A1(n20277), .O(n20666) );
  INV2 U22630 ( .I(n20666), .O(n21093) );
  XNR2HS U22631 ( .I1(n20872), .I2(n21393), .O(n20280) );
  XNR2HS U22632 ( .I1(n20280), .I2(n21472), .O(n20664) );
  INV1S U22633 ( .I(n20664), .O(n20642) );
  AOI22S U22634 ( .A1(n20286), .A2(n20364), .B1(n20363), .B2(n20286), .O(
        n20290) );
  ND2S U22635 ( .I1(n20281), .I2(n19818), .O(n20284) );
  ND2S U22636 ( .I1(n21259), .I2(n18142), .O(n20282) );
  ND2S U22637 ( .I1(n20287), .I2(n20373), .O(n20288) );
  INV1S U22638 ( .I(n20291), .O(n20292) );
  MXL2H U22639 ( .A(n22661), .B(n20292), .S(n13822), .OB(n23845) );
  INV1S U22640 ( .I(n29503), .O(n20313) );
  AOI22S U22641 ( .A1(n20298), .A2(n20371), .B1(n20364), .B2(n20298), .O(
        n20302) );
  ND2S U22642 ( .I1(n21254), .I2(n18142), .O(n20294) );
  ND2S U22643 ( .I1(n20299), .I2(n20373), .O(n20300) );
  OR2P U22644 ( .I1(n13822), .I2(n22662), .O(n21191) );
  OAI12HP U22645 ( .B1(n20809), .B2(n20685), .A1(n21191), .O(n24768) );
  AOI22S U22646 ( .A1(n20308), .A2(n20363), .B1(n20364), .B2(n20308), .O(
        n20312) );
  ND2S U22647 ( .I1(n20303), .I2(n19818), .O(n20306) );
  ND2S U22648 ( .I1(n20366), .I2(n20303), .O(n20305) );
  ND2S U22649 ( .I1(n21245), .I2(n18142), .O(n20304) );
  AOI12HS U22650 ( .B1(n20308), .B2(n20371), .A1(n20307), .O(n20311) );
  ND2S U22651 ( .I1(n20309), .I2(n20373), .O(n20310) );
  MXL2HP U22652 ( .A(n22663), .B(n20688), .S(n13822), .OB(n26012) );
  MOAI1S U22653 ( .A1(n20313), .A2(n24768), .B1(n21596), .B2(n21595), .O(
        n20381) );
  AOI22S U22654 ( .A1(n20320), .A2(n20363), .B1(n20314), .B2(n20320), .O(
        n20323) );
  ND2S U22655 ( .I1(n20315), .I2(n19818), .O(n20318) );
  ND2S U22656 ( .I1(n20366), .I2(n20315), .O(n20317) );
  ND2S U22657 ( .I1(n22932), .I2(n18142), .O(n20316) );
  ND3S U22658 ( .I1(n20318), .I2(n20317), .I3(n20316), .O(n20319) );
  AOI12HS U22659 ( .B1(n20320), .B2(n20364), .A1(n20319), .O(n20322) );
  ND3HT U22660 ( .I1(n20323), .I2(n20322), .I3(n20321), .O(n22671) );
  ND2S U22661 ( .I1(n20324), .I2(n19818), .O(n20327) );
  ND2S U22662 ( .I1(n20366), .I2(n20324), .O(n20326) );
  ND2S U22663 ( .I1(n13887), .I2(n18142), .O(n20325) );
  ND3 U22664 ( .I1(n20327), .I2(n20326), .I3(n20325), .O(n20328) );
  AOI12HS U22665 ( .B1(n20329), .B2(n20371), .A1(n20328), .O(n20333) );
  AOI22S U22666 ( .A1(n20329), .A2(n20364), .B1(n20363), .B2(n20329), .O(
        n20332) );
  ND2S U22667 ( .I1(n20330), .I2(n20373), .O(n20331) );
  ND3HT U22668 ( .I1(n20333), .I2(n20332), .I3(n20331), .O(n22668) );
  AOI22S U22669 ( .A1(n20339), .A2(n20371), .B1(n20363), .B2(n20339), .O(
        n20342) );
  ND2S U22670 ( .I1(n20334), .I2(n19818), .O(n20337) );
  ND2S U22671 ( .I1(n20366), .I2(n20334), .O(n20336) );
  ND2S U22672 ( .I1(n21225), .I2(n18142), .O(n20335) );
  AOI12HS U22673 ( .B1(n20339), .B2(n20364), .A1(n20338), .O(n20341) );
  ND3P U22674 ( .I1(n20342), .I2(n20341), .I3(n20340), .O(n22667) );
  ND2S U22675 ( .I1(n20644), .I2(n22713), .O(n20356) );
  MXL2HP U22676 ( .A(n22668), .B(n20343), .S(n13822), .OB(n26638) );
  ND2S U22677 ( .I1(n20344), .I2(n19818), .O(n20348) );
  ND2S U22678 ( .I1(n20366), .I2(n20344), .O(n20347) );
  ND2S U22679 ( .I1(n20351), .I2(n20373), .O(n20352) );
  ND3HT U22680 ( .I1(n20354), .I2(n20353), .I3(n20352), .O(n22670) );
  INV1S U22681 ( .I(n22670), .O(n20810) );
  OAI112HS U22682 ( .C1(n26638), .C2(n21810), .A1(n21635), .B1(n20810), .O(
        n20355) );
  OAI112HS U22683 ( .C1(n29461), .C2(n22668), .A1(n20356), .B1(n20355), .O(
        n20361) );
  MXL2HP U22684 ( .A(n22671), .B(n20357), .S(n13822), .OB(n27262) );
  INV2 U22685 ( .I(n27262), .O(n29444) );
  ND2S U22686 ( .I1(n29442), .I2(n29444), .O(n20360) );
  INV2 U22687 ( .I(n25391), .O(n29485) );
  ND2S U22688 ( .I1(n29483), .I2(n29485), .O(n20359) );
  ND3 U22689 ( .I1(n20361), .I2(n20360), .I3(n20359), .O(n20362) );
  OAI12HS U22690 ( .B1(n29442), .B2(n22671), .A1(n20362), .O(n20379) );
  ND2S U22691 ( .I1(n20365), .I2(n19818), .O(n20369) );
  ND2S U22692 ( .I1(n20366), .I2(n20365), .O(n20368) );
  ND3 U22693 ( .I1(n20369), .I2(n20368), .I3(n20367), .O(n20370) );
  AOI12HS U22694 ( .B1(n20372), .B2(n20371), .A1(n20370), .O(n20376) );
  ND2S U22695 ( .I1(n20374), .I2(n20373), .O(n20375) );
  MXL2HP U22696 ( .A(n22669), .B(n21655), .S(n13822), .OB(n28528) );
  NR2 U22697 ( .I1(n22663), .I2(n21595), .O(n20378) );
  AOI12HS U22698 ( .B1(n20379), .B2(n13938), .A1(n13937), .O(n20380) );
  OAI22S U22699 ( .A1(n20381), .A2(n20380), .B1(n22662), .B2(n29503), .O(
        n20382) );
  OAI12HS U22700 ( .B1(n23845), .B2(n20383), .A1(n20382), .O(n20384) );
  OAI12HS U22701 ( .B1(n21467), .B2(n22661), .A1(n20384), .O(n21194) );
  NR2 U22702 ( .I1(n21653), .I2(n29503), .O(n20401) );
  MXL2H U22703 ( .A(n29448), .B(n20679), .S(n21654), .OB(n29441) );
  OAI22S U22704 ( .A1(n21611), .A2(n20740), .B1(n29442), .B2(n29441), .O(
        n20395) );
  ND2P U22705 ( .I1(n13887), .I2(n20809), .O(n29467) );
  ND2S U22706 ( .I1(n29461), .I2(n21658), .O(n20387) );
  INV1S U22707 ( .I(n21657), .O(n20735) );
  ND3S U22708 ( .I1(n20387), .I2(n21635), .I3(n20735), .O(n20393) );
  ND2S U22709 ( .I1(n20643), .I2(n22331), .O(n20392) );
  NR2T U22710 ( .I1(n13822), .I2(n13818), .O(n21246) );
  NR2 U22711 ( .I1(n21246), .I2(n21654), .O(n20389) );
  AN2 U22712 ( .I1(n20388), .I2(n21654), .O(n20678) );
  NR2T U22713 ( .I1(n20389), .I2(n20678), .O(n21659) );
  ND2S U22714 ( .I1(n20644), .I2(n13813), .O(n20391) );
  ND2T U22715 ( .I1(n21659), .I2(n20809), .O(n20769) );
  OAI22S U22716 ( .A1(n13815), .A2(n21811), .B1(n21812), .B2(n20769), .O(
        n20390) );
  AOI13HS U22717 ( .B1(n20393), .B2(n20392), .B3(n20391), .A1(n20390), .O(
        n20394) );
  OR2 U22718 ( .I1(n13822), .I2(n20757), .O(n20776) );
  OAI22S U22719 ( .A1(n20395), .A2(n20394), .B1(n21808), .B2(n20776), .O(
        n20399) );
  ND2P U22720 ( .I1(n21660), .I2(n20809), .O(n20780) );
  OAI22S U22721 ( .A1(n20780), .A2(n21805), .B1(n21804), .B2(n20784), .O(
        n20397) );
  AOI12HS U22722 ( .B1(n20399), .B2(n20398), .A1(n20397), .O(n20400) );
  OAI22S U22723 ( .A1(n20401), .A2(n20400), .B1(n20788), .B2(n21803), .O(
        n20402) );
  OAI12HS U22724 ( .B1(n21669), .B2(n21467), .A1(n20402), .O(n20796) );
  INV1S U22725 ( .I(n20796), .O(n20792) );
  INV1S U22726 ( .I(n20403), .O(n20405) );
  MOAI1S U22727 ( .A1(n13929), .A2(n20405), .B1(n20404), .B2(n20438), .O(
        n20410) );
  MOAI1S U22728 ( .A1(n13946), .A2(n20408), .B1(n20407), .B2(n20406), .O(
        n20409) );
  NR2 U22729 ( .I1(n20410), .I2(n20409), .O(n20417) );
  AOI22S U22730 ( .A1(n20412), .A2(n13846), .B1(n13839), .B2(n20411), .O(
        n20416) );
  AOI22S U22731 ( .A1(n20414), .A2(n13791), .B1(n20963), .B2(n20413), .O(
        n20415) );
  ND3S U22732 ( .I1(n20417), .I2(n20416), .I3(n20415), .O(n20434) );
  INV1S U22733 ( .I(n20418), .O(n20420) );
  MOAI1S U22734 ( .A1(n20421), .A2(n20420), .B1(n20419), .B2(n17762), .O(
        n20425) );
  MOAI1S U22735 ( .A1(n13844), .A2(n20423), .B1(n20422), .B2(n17928), .O(
        n20424) );
  NR2 U22736 ( .I1(n20425), .I2(n20424), .O(n20432) );
  AOI22S U22737 ( .A1(n20427), .A2(n17875), .B1(n20613), .B2(n20426), .O(
        n20431) );
  AOI22S U22738 ( .A1(n20429), .A2(n21062), .B1(n13830), .B2(n20428), .O(
        n20430) );
  ND3S U22739 ( .I1(n20432), .I2(n20431), .I3(n20430), .O(n20433) );
  NR2 U22740 ( .I1(n20434), .I2(n20433), .O(n20435) );
  ND2S U22741 ( .I1(n21812), .I2(n21330), .O(n20506) );
  NR2P U22742 ( .I1(n13822), .I2(n21221), .O(n21329) );
  ND2S U22743 ( .I1(n21809), .I2(n21329), .O(n20467) );
  AOI22S U22744 ( .A1(n20440), .A2(n20439), .B1(n20438), .B2(n20437), .O(
        n20450) );
  AOI22S U22745 ( .A1(n20442), .A2(n19914), .B1(n13847), .B2(n20441), .O(
        n20449) );
  AOI22S U22746 ( .A1(n20444), .A2(n13846), .B1(n13839), .B2(n20443), .O(
        n20448) );
  AOI22S U22747 ( .A1(n20446), .A2(n13791), .B1(n20187), .B2(n20445), .O(
        n20447) );
  AN4S U22748 ( .I1(n20450), .I2(n20449), .I3(n20448), .I4(n20447), .O(n20464)
         );
  AOI22S U22749 ( .A1(n20452), .A2(n20613), .B1(n17875), .B2(n20451), .O(
        n20462) );
  AOI22S U22750 ( .A1(n20454), .A2(n21062), .B1(n13830), .B2(n20453), .O(
        n20461) );
  AOI22S U22751 ( .A1(n20456), .A2(n17762), .B1(n20560), .B2(n20455), .O(
        n20460) );
  AOI22S U22752 ( .A1(n20458), .A2(n20969), .B1(n17928), .B2(n20457), .O(
        n20459) );
  AN4S U22753 ( .I1(n20462), .I2(n20461), .I3(n20460), .I4(n20459), .O(n20463)
         );
  ND2S U22754 ( .I1(n20464), .I2(n20463), .O(n20465) );
  NR2 U22755 ( .I1(n26639), .I2(n20643), .O(n20466) );
  OAI22S U22756 ( .A1(n20467), .A2(n20466), .B1(n29461), .B2(n21333), .O(
        n20501) );
  AOI22S U22757 ( .A1(n20469), .A2(n13835), .B1(n20263), .B2(n20468), .O(
        n20473) );
  AOI22S U22758 ( .A1(n20471), .A2(n13839), .B1(n13847), .B2(n20470), .O(
        n20472) );
  ND2S U22759 ( .I1(n20473), .I2(n20472), .O(n20498) );
  AOI22S U22760 ( .A1(n20475), .A2(n13846), .B1(n20963), .B2(n20474), .O(
        n20479) );
  AOI22S U22761 ( .A1(n20477), .A2(n20613), .B1(n13791), .B2(n20476), .O(
        n20478) );
  ND2S U22762 ( .I1(n20479), .I2(n20478), .O(n20497) );
  ND2S U22763 ( .I1(n20480), .I2(n17928), .O(n20483) );
  ND2S U22764 ( .I1(n20481), .I2(n20620), .O(n20482) );
  ND3S U22765 ( .I1(n20483), .I2(n20482), .I3(n13822), .O(n20488) );
  INV1S U22766 ( .I(n20484), .O(n20486) );
  MOAI1S U22767 ( .A1(n13844), .A2(n20486), .B1(n20485), .B2(n17762), .O(
        n20487) );
  NR2 U22768 ( .I1(n20488), .I2(n20487), .O(n20495) );
  AOI22S U22769 ( .A1(n20490), .A2(n13830), .B1(n17875), .B2(n20489), .O(
        n20494) );
  AOI22S U22770 ( .A1(n20492), .A2(n21062), .B1(n21061), .B2(n20491), .O(
        n20493) );
  ND3S U22771 ( .I1(n20495), .I2(n20494), .I3(n20493), .O(n20496) );
  NR3 U22772 ( .I1(n20498), .I2(n20497), .I3(n20496), .O(n20499) );
  AOI22S U22773 ( .A1(n29445), .A2(n29442), .B1(n29483), .B2(n29486), .O(
        n20500) );
  ND2 U22774 ( .I1(n20501), .I2(n20500), .O(n20505) );
  ND2S U22775 ( .I1(n20506), .I2(n21228), .O(n20502) );
  ND2S U22776 ( .I1(n20503), .I2(n20502), .O(n20504) );
  OAI112HS U22777 ( .C1(n29445), .C2(n20506), .A1(n20505), .B1(n20504), .O(
        n20536) );
  AOI22S U22778 ( .A1(n20508), .A2(n20263), .B1(n20438), .B2(n20507), .O(
        n20518) );
  AOI22S U22779 ( .A1(n20510), .A2(n19914), .B1(n13847), .B2(n20509), .O(
        n20517) );
  AOI22S U22780 ( .A1(n20512), .A2(n13846), .B1(n13839), .B2(n20511), .O(
        n20516) );
  AOI22S U22781 ( .A1(n20514), .A2(n13791), .B1(n20187), .B2(n20513), .O(
        n20515) );
  AN4S U22782 ( .I1(n20518), .I2(n20517), .I3(n20516), .I4(n20515), .O(n20533)
         );
  AOI22S U22783 ( .A1(n20520), .A2(n20613), .B1(n17875), .B2(n20519), .O(
        n20531) );
  AOI22S U22784 ( .A1(n20522), .A2(n19483), .B1(n13830), .B2(n20521), .O(
        n20530) );
  AOI22S U22785 ( .A1(n20525), .A2(n17762), .B1(n20524), .B2(n20523), .O(
        n20529) );
  AOI22S U22786 ( .A1(n20527), .A2(n20969), .B1(n17928), .B2(n20526), .O(
        n20528) );
  AN4S U22787 ( .I1(n20531), .I2(n20530), .I3(n20529), .I4(n20528), .O(n20532)
         );
  ND2S U22788 ( .I1(n20533), .I2(n20532), .O(n20534) );
  MXL2H U22789 ( .A(n20534), .B(n20711), .S(n20809), .OB(n28531) );
  MAO222 U22790 ( .A1(n20536), .B1(n28531), .C1(n20535), .O(n20604) );
  INV1S U22791 ( .I(n21340), .O(n20538) );
  NR2 U22792 ( .I1(n20538), .I2(n13814), .O(n20603) );
  AOI22S U22793 ( .A1(n20540), .A2(n13793), .B1(n20263), .B2(n20539), .O(
        n20550) );
  AOI22S U22794 ( .A1(n20542), .A2(n13839), .B1(n13847), .B2(n20541), .O(
        n20549) );
  AOI22S U22795 ( .A1(n20544), .A2(n13846), .B1(n20963), .B2(n20543), .O(
        n20548) );
  AOI22S U22796 ( .A1(n20546), .A2(n13791), .B1(n20613), .B2(n20545), .O(
        n20547) );
  AN4S U22797 ( .I1(n20550), .I2(n20549), .I3(n20548), .I4(n20547), .O(n20568)
         );
  ND2S U22798 ( .I1(n20551), .I2(n17928), .O(n20554) );
  ND2S U22799 ( .I1(n20552), .I2(n20620), .O(n20553) );
  ND3S U22800 ( .I1(n20554), .I2(n20553), .I3(n13822), .O(n20566) );
  MOAI1S U22801 ( .A1(n13844), .A2(n20556), .B1(n20555), .B2(n17762), .O(
        n20565) );
  AOI22S U22802 ( .A1(n20558), .A2(n13830), .B1(n17875), .B2(n20557), .O(
        n20563) );
  AOI22S U22803 ( .A1(n20561), .A2(n19483), .B1(n20560), .B2(n20559), .O(
        n20562) );
  NR3 U22804 ( .I1(n20566), .I2(n20565), .I3(n20564), .O(n20567) );
  ND2S U22805 ( .I1(n20569), .I2(n17928), .O(n20572) );
  ND2S U22806 ( .I1(n20570), .I2(n20620), .O(n20571) );
  MOAI1S U22807 ( .A1(n13844), .A2(n20574), .B1(n20573), .B2(n17762), .O(
        n20575) );
  NR2 U22808 ( .I1(n20576), .I2(n20575), .O(n20584) );
  AOI22S U22809 ( .A1(n20578), .A2(n13830), .B1(n17875), .B2(n20577), .O(
        n20583) );
  AOI22S U22810 ( .A1(n20581), .A2(n21062), .B1(n20580), .B2(n20579), .O(
        n20582) );
  MOAI1S U22811 ( .A1(n13946), .A2(n20589), .B1(n20588), .B2(n13839), .O(
        n20590) );
  NR2 U22812 ( .I1(n20591), .I2(n20590), .O(n20598) );
  AOI22S U22813 ( .A1(n20593), .A2(n13846), .B1(n14174), .B2(n20592), .O(
        n20597) );
  AOI22S U22814 ( .A1(n20595), .A2(n13791), .B1(n20613), .B2(n20594), .O(
        n20596) );
  ND3S U22815 ( .I1(n20598), .I2(n20597), .I3(n20596), .O(n20599) );
  NR2 U22816 ( .I1(n20600), .I2(n20599), .O(n20601) );
  AOI22S U22817 ( .A1(n21595), .A2(n21597), .B1(n29509), .B2(n29503), .O(
        n20602) );
  OA12P U22818 ( .B1(n20604), .B2(n20603), .A1(n20602), .O(n20639) );
  NR2 U22819 ( .I1(n20605), .I2(n29503), .O(n20638) );
  AOI22S U22820 ( .A1(n20607), .A2(n19914), .B1(n20439), .B2(n20606), .O(
        n20618) );
  AOI22S U22821 ( .A1(n20609), .A2(n13839), .B1(n13847), .B2(n20608), .O(
        n20617) );
  AOI22S U22822 ( .A1(n20611), .A2(n13846), .B1(n20187), .B2(n20610), .O(
        n20616) );
  AOI22S U22823 ( .A1(n20614), .A2(n13791), .B1(n20613), .B2(n20612), .O(
        n20615) );
  AN4S U22824 ( .I1(n20618), .I2(n20617), .I3(n20616), .I4(n20615), .O(n20637)
         );
  ND2S U22825 ( .I1(n20619), .I2(n17928), .O(n20623) );
  ND2S U22826 ( .I1(n20621), .I2(n20620), .O(n20622) );
  ND3S U22827 ( .I1(n20623), .I2(n20622), .I3(n13822), .O(n20635) );
  MOAI1S U22828 ( .A1(n13844), .A2(n20625), .B1(n20624), .B2(n17762), .O(
        n20634) );
  AOI22S U22829 ( .A1(n20627), .A2(n13830), .B1(n17875), .B2(n20626), .O(
        n20632) );
  AOI22S U22830 ( .A1(n20630), .A2(n21062), .B1(n20629), .B2(n20628), .O(
        n20631) );
  NR3 U22831 ( .I1(n20635), .I2(n20634), .I3(n20633), .O(n20636) );
  MOAI1H U22832 ( .A1(n20639), .A2(n20638), .B1(n21460), .B2(n21467), .O(
        n20640) );
  XOR2HS U22833 ( .I1(n20792), .I2(n21353), .O(n20641) );
  XNR2HS U22834 ( .I1(n21206), .I2(n20641), .O(n20665) );
  ND2S U22835 ( .I1(n20642), .I2(n20665), .O(n20660) );
  AOI12HS U22836 ( .B1(n20662), .B2(n21093), .A1(n20660), .O(n20661) );
  ND2S U22837 ( .I1(n20643), .I2(n15985), .O(n20648) );
  ND2S U22838 ( .I1(n20644), .I2(n13818), .O(n20647) );
  OAI112HS U22839 ( .C1(n15985), .C2(n21810), .A1(n21635), .B1(n22942), .O(
        n20646) );
  INV1S U22840 ( .I(n21246), .O(n29489) );
  MOAI1S U22841 ( .A1(n20644), .A2(n29489), .B1(n21117), .B2(n21910), .O(
        n20645) );
  AOI13HS U22842 ( .B1(n20648), .B2(n20647), .B3(n20646), .A1(n20645), .O(
        n20650) );
  OAI22S U22843 ( .A1(n20863), .A2(n21611), .B1(n29442), .B2(n22932), .O(
        n20649) );
  ND2P U22844 ( .I1(n20863), .I2(n20809), .O(n21616) );
  OAI22S U22845 ( .A1(n20650), .A2(n20649), .B1(n21808), .B2(n21616), .O(
        n20651) );
  OR2 U22846 ( .I1(n29513), .I2(n21804), .O(n20652) );
  ND2S U22847 ( .I1(n21280), .I2(n20666), .O(n20657) );
  MAO222 U22848 ( .A1(n20796), .B1(n21353), .C1(n21194), .O(n20656) );
  XOR2HS U22849 ( .I1(n20657), .I2(n20656), .O(n20658) );
  XNR2HS U22850 ( .I1(n20658), .I2(n20662), .O(n20663) );
  INV1S U22851 ( .I(n20663), .O(n20659) );
  MXL2HS U22852 ( .A(n20661), .B(n20660), .S(n20659), .OB(n20673) );
  OAI12HS U22853 ( .B1(n20663), .B2(n20662), .A1(n20666), .O(n20667) );
  XNR2HS U22854 ( .I1(n20665), .I2(n20664), .O(n20668) );
  MXL2HS U22855 ( .A(n20667), .B(n20666), .S(n20668), .OB(n20671) );
  XNR2HS U22856 ( .I1(n21093), .I2(n20669), .O(n20670) );
  INV1S U22857 ( .I(n21280), .O(n21283) );
  MXL2HS U22858 ( .A(n20671), .B(n20670), .S(n21283), .OB(n20672) );
  ND2P U22859 ( .I1(n21658), .I2(n20809), .O(n20765) );
  OR2 U22860 ( .I1(n21225), .I2(n20769), .O(n20677) );
  AN2 U22861 ( .I1(n21657), .I2(n20809), .O(n21644) );
  ND2S U22862 ( .I1(n20674), .I2(n13887), .O(n20675) );
  ND3S U22863 ( .I1(n21644), .I2(n22942), .I3(n20675), .O(n20676) );
  OAI112HS U22864 ( .C1(n20765), .C2(n13887), .A1(n20677), .B1(n20676), .O(
        n20682) );
  AOI22S U22865 ( .A1(n20679), .A2(n21117), .B1(n20678), .B2(n21246), .O(
        n20681) );
  MOAI1S U22866 ( .A1(n20776), .A2(n20863), .B1(n13816), .B2(n29441), .O(
        n20680) );
  AOI12HS U22867 ( .B1(n20682), .B2(n20681), .A1(n20680), .O(n20684) );
  NR2 U22868 ( .I1(n21616), .I2(n20740), .O(n20683) );
  INV1S U22869 ( .I(n20780), .O(n21594) );
  MOAI1S U22870 ( .A1(n20684), .A2(n20683), .B1(n23508), .B2(n21594), .O(
        n20687) );
  OR2S U22871 ( .I1(n20685), .I2(n29513), .O(n20686) );
  OAI112HS U22872 ( .C1(n19494), .C2(n20688), .A1(n20687), .B1(n20686), .O(
        n20690) );
  AOI22S U22873 ( .A1(n20691), .A2(n21237), .B1(n20690), .B2(n20689), .O(
        n21286) );
  INV1S U22874 ( .I(n21286), .O(n21220) );
  INV1S U22875 ( .I(n20788), .O(n21392) );
  INV1S U22876 ( .I(n20776), .O(n21610) );
  OR2 U22877 ( .I1(n21658), .I2(n21072), .O(n20693) );
  OAI22S U22878 ( .A1(n20769), .A2(n23186), .B1(n23188), .B2(n20765), .O(
        n20692) );
  AOI13HS U22879 ( .B1(n20693), .B2(n21644), .B3(n23427), .A1(n20692), .O(
        n20694) );
  OAI22S U22880 ( .A1(n20695), .A2(n20694), .B1(n13815), .B2(n20942), .O(
        n20696) );
  OAI12HS U22881 ( .B1(n21610), .B2(n21023), .A1(n20696), .O(n20699) );
  INV1S U22882 ( .I(n20784), .O(n29501) );
  OAI22S U22883 ( .A1(n29501), .A2(n21088), .B1(n21081), .B2(n21594), .O(
        n20697) );
  AO12 U22884 ( .B1(n20699), .B2(n20698), .A1(n20697), .O(n20702) );
  OAI12HS U22885 ( .B1(n21392), .B2(n21085), .A1(n20703), .O(n21090) );
  OR2 U22886 ( .I1(n21220), .I2(n21090), .O(n20804) );
  INV1S U22887 ( .I(n20804), .O(n20705) );
  INV1S U22888 ( .I(n21090), .O(n21096) );
  NR2 U22889 ( .I1(n21286), .I2(n21096), .O(n20704) );
  NR2 U22890 ( .I1(n20705), .I2(n20704), .O(n20750) );
  ND2S U22891 ( .I1(n29441), .I2(n20809), .O(n20722) );
  ND2S U22892 ( .I1(n21657), .I2(n21329), .O(n20707) );
  NR2 U22893 ( .I1(n21658), .I2(n26639), .O(n20706) );
  NR2 U22894 ( .I1(n20707), .I2(n20706), .O(n20709) );
  MOAI1S U22895 ( .A1(n20765), .A2(n21333), .B1(n21659), .B2(n21330), .O(
        n20708) );
  MOAI1S U22896 ( .A1(n20709), .A2(n20708), .B1(n29486), .B2(n20769), .O(
        n20710) );
  OAI12HS U22897 ( .B1(n21228), .B2(n20722), .A1(n20710), .O(n20714) );
  INV1S U22898 ( .I(n28531), .O(n21613) );
  AOI22S U22899 ( .A1(n29445), .A2(n13815), .B1(n21613), .B2(n20776), .O(
        n20713) );
  MOAI1S U22900 ( .A1(n20776), .A2(n20711), .B1(n21340), .B2(n21660), .O(
        n20712) );
  AOI12HS U22901 ( .B1(n20714), .B2(n20713), .A1(n20712), .O(n20716) );
  MOAI1S U22902 ( .A1(n21594), .A2(n26013), .B1(n29509), .B2(n20784), .O(
        n20715) );
  MOAI1S U22903 ( .A1(n20716), .A2(n20715), .B1(n21345), .B2(n21653), .O(
        n20717) );
  OAI12HS U22904 ( .B1(n21392), .B2(n23846), .A1(n20717), .O(n20718) );
  OAI12HS U22905 ( .B1(n21236), .B2(n20788), .A1(n20718), .O(n21350) );
  INV1S U22906 ( .I(n20765), .O(n29460) );
  OR2 U22907 ( .I1(n29460), .I2(n26638), .O(n20721) );
  INV1S U22908 ( .I(n21644), .O(n20719) );
  OAI22S U22909 ( .A1(n20765), .A2(n22668), .B1(n22670), .B2(n20719), .O(
        n20720) );
  OAI112HS U22910 ( .C1(n25391), .C2(n29493), .A1(n20721), .B1(n20720), .O(
        n20724) );
  OR2 U22911 ( .I1(n20722), .I2(n22671), .O(n20723) );
  OAI112HS U22912 ( .C1(n22667), .C2(n20769), .A1(n20724), .B1(n20723), .O(
        n20727) );
  ND3S U22913 ( .I1(n20727), .I2(n20726), .I3(n20725), .O(n20731) );
  INV1S U22914 ( .I(n22663), .O(n20728) );
  AOI22S U22915 ( .A1(n21594), .A2(n20728), .B1(n28528), .B2(n21610), .O(
        n20730) );
  OAI22S U22916 ( .A1(n29501), .A2(n24768), .B1(n26012), .B2(n21594), .O(
        n20729) );
  AOI12HS U22917 ( .B1(n20731), .B2(n20730), .A1(n20729), .O(n20734) );
  OAI22S U22918 ( .A1(n22302), .A2(n21191), .B1(n22661), .B2(n20788), .O(
        n20733) );
  OA12 U22919 ( .B1(n20734), .B2(n20733), .A1(n20732), .O(n21154) );
  INV1S U22920 ( .I(n21154), .O(n21203) );
  XOR2HS U22921 ( .I1(n21350), .I2(n21203), .O(n20749) );
  OAI22S U22922 ( .A1(n20780), .A2(n22412), .B1(n22411), .B2(n20784), .O(
        n20746) );
  INV1S U22923 ( .I(n20903), .O(n21602) );
  ND2T U22924 ( .I1(n22417), .I2(n20809), .O(n29470) );
  OAI112HS U22925 ( .C1(n22417), .C2(n22331), .A1(n20735), .B1(n22419), .O(
        n20736) );
  OAI112HS U22926 ( .C1(n20891), .C2(n21659), .A1(n20737), .B1(n20736), .O(
        n20739) );
  OA22 U22927 ( .A1(n13815), .A2(n22415), .B1(n22416), .B2(n20769), .O(n20738)
         );
  ND2S U22928 ( .I1(n20739), .I2(n20738), .O(n20742) );
  ND2S U22929 ( .I1(n20742), .I2(n20741), .O(n20744) );
  AOI22S U22930 ( .A1(n22322), .A2(n21602), .B1(n20744), .B2(n20743), .O(
        n20745) );
  OAI22S U22931 ( .A1(n20746), .A2(n20745), .B1(n21653), .B2(n29519), .O(
        n20748) );
  AOI22S U22932 ( .A1(n21391), .A2(n22324), .B1(n20748), .B2(n20747), .O(
        n20921) );
  XNR2HS U22933 ( .I1(n20749), .I2(n20840), .O(n20795) );
  XOR2HS U22934 ( .I1(n20750), .I2(n20795), .O(n20794) );
  NR2 U22935 ( .I1(n20776), .I2(n22062), .O(n20759) );
  INV2 U22936 ( .I(n21407), .O(n21618) );
  AN2S U22937 ( .I1(n21399), .I2(n29493), .O(n20754) );
  INV1S U22938 ( .I(n21643), .O(n21177) );
  OAI22S U22939 ( .A1(n21658), .A2(n21394), .B1(n21177), .B2(n21657), .O(
        n20752) );
  ND2S U22940 ( .I1(n21394), .I2(n21658), .O(n20751) );
  AOI22S U22941 ( .A1(n29491), .A2(n13813), .B1(n20752), .B2(n20751), .O(
        n20753) );
  OAI22S U22942 ( .A1(n20754), .A2(n20753), .B1(n29441), .B2(n21403), .O(
        n20756) );
  OR2S U22943 ( .I1(n13815), .I2(n22059), .O(n20755) );
  AOI22S U22944 ( .A1(n20757), .A2(n21618), .B1(n20756), .B2(n20755), .O(
        n20758) );
  OAI22S U22945 ( .A1(n20759), .A2(n20758), .B1(n21660), .B2(n21412), .O(
        n20761) );
  OAI112HS U22946 ( .C1(n22055), .C2(n20780), .A1(n20761), .B1(n20760), .O(
        n20763) );
  AOI22H U22947 ( .A1(n21392), .A2(n13809), .B1(n20763), .B2(n20762), .O(
        n21435) );
  NR2 U22948 ( .I1(n20769), .I2(n29497), .O(n20764) );
  NR2 U22949 ( .I1(n13815), .I2(n29455), .O(n20772) );
  NR2 U22950 ( .I1(n20764), .I2(n20772), .O(n20775) );
  NR2 U22951 ( .I1(n20765), .I2(n29475), .O(n20768) );
  AN2S U22952 ( .I1(n27893), .I2(n21644), .O(n20767) );
  ND2S U22953 ( .I1(n29475), .I2(n20765), .O(n20766) );
  OAI12HS U22954 ( .B1(n20768), .B2(n20767), .A1(n20766), .O(n20774) );
  ND2S U22955 ( .I1(n29497), .I2(n20769), .O(n20771) );
  ND2S U22956 ( .I1(n29455), .I2(n13815), .O(n20770) );
  OAI12HS U22957 ( .B1(n20772), .B2(n20771), .A1(n20770), .O(n20773) );
  AOI12HS U22958 ( .B1(n20775), .B2(n20774), .A1(n20773), .O(n20779) );
  NR2 U22959 ( .I1(n20776), .I2(n28527), .O(n20778) );
  ND2S U22960 ( .I1(n28527), .I2(n20776), .O(n20777) );
  OAI12HS U22961 ( .B1(n20779), .B2(n20778), .A1(n20777), .O(n20783) );
  OR2 U22962 ( .I1(n20780), .I2(n21411), .O(n20782) );
  AOI12HS U22963 ( .B1(n20783), .B2(n20782), .A1(n20781), .O(n20787) );
  NR2 U22964 ( .I1(n20784), .I2(n21416), .O(n20786) );
  OAI12HS U22965 ( .B1(n20787), .B2(n20786), .A1(n20785), .O(n20791) );
  OR2 U22966 ( .I1(n20788), .I2(n23839), .O(n20790) );
  XOR2HS U22967 ( .I1(n20792), .I2(n13909), .O(n20793) );
  XNR2HS U22968 ( .I1(n21435), .I2(n20793), .O(n20801) );
  INV1S U22969 ( .I(n20801), .O(n20800) );
  XNR2HS U22970 ( .I1(n20794), .I2(n20800), .O(n20808) );
  ND2S U22971 ( .I1(n20795), .I2(n20804), .O(n20799) );
  NR2 U22972 ( .I1(n20796), .I2(n13909), .O(n20798) );
  MOAI1S U22973 ( .A1(n20798), .A2(n20797), .B1(n13909), .B2(n20796), .O(
        n20803) );
  INV1S U22974 ( .I(n21350), .O(n21356) );
  MAO222 U22975 ( .A1(n20840), .B1(n21356), .C1(n21203), .O(n20802) );
  MOAI1 U22976 ( .A1(n20800), .A2(n20799), .B1(n20803), .B2(n20802), .O(n20806) );
  OAI22S U22977 ( .A1(n20801), .A2(n20804), .B1(n20803), .B2(n20802), .O(
        n20805) );
  XOR2HS U22978 ( .I1(n20806), .I2(n20805), .O(n20807) );
  INV2 U22979 ( .I(n24768), .O(n29508) );
  INV1 U22980 ( .I(n28528), .O(n21612) );
  INV2 U22981 ( .I(n26638), .O(n29463) );
  ND3S U22982 ( .I1(n22419), .I2(n20810), .I3(n20809), .O(n20811) );
  OR2 U22983 ( .I1(n22667), .I2(n20891), .O(n20812) );
  ND3 U22984 ( .I1(n20814), .I2(n20813), .I3(n20812), .O(n20817) );
  ND2S U22985 ( .I1(n20891), .I2(n29485), .O(n20816) );
  ND2S U22986 ( .I1(n20892), .I2(n29444), .O(n20815) );
  ND3P U22987 ( .I1(n20817), .I2(n20816), .I3(n20815), .O(n20819) );
  NR2 U22988 ( .I1(n21612), .I2(n20899), .O(n20820) );
  OR2 U22989 ( .I1(n22663), .I2(n20903), .O(n20822) );
  AOI22H U22990 ( .A1(n29508), .A2(n29519), .B1(n20823), .B2(n20822), .O(
        n20825) );
  NR2 U22991 ( .I1(n21191), .I2(n13811), .O(n20824) );
  INV1S U22992 ( .I(n23845), .O(n21457) );
  MOAI1H U22993 ( .A1(n20825), .A2(n20824), .B1(n21457), .B2(n19461), .O(
        n20826) );
  ND2S U22994 ( .I1(n22419), .I2(n21329), .O(n20828) );
  NR2 U22995 ( .I1(n26639), .I2(n22417), .O(n20827) );
  MAOI1 U22996 ( .A1(n21330), .A2(n22416), .B1(n20828), .B2(n20827), .O(n20829) );
  OAI12HS U22997 ( .B1(n29470), .B2(n21333), .A1(n20829), .O(n20832) );
  ND2S U22998 ( .I1(n20891), .I2(n29486), .O(n20831) );
  ND2S U22999 ( .I1(n20892), .I2(n29445), .O(n20830) );
  ND3 U23000 ( .I1(n20832), .I2(n20831), .I3(n20830), .O(n20833) );
  OAI12HS U23001 ( .B1(n21228), .B2(n20892), .A1(n20833), .O(n20834) );
  INV1S U23002 ( .I(n20899), .O(n21619) );
  MAO222 U23003 ( .A1(n20834), .B1(n28531), .C1(n21619), .O(n20837) );
  AOI22S U23004 ( .A1(n29519), .A2(n29509), .B1(n21597), .B2(n20903), .O(
        n20835) );
  OAI12HS U23005 ( .B1(n20837), .B2(n20836), .A1(n20835), .O(n20839) );
  AOI22S U23006 ( .A1(n22410), .A2(n21346), .B1(n21345), .B2(n22411), .O(
        n20838) );
  AOI22S U23007 ( .A1(n21460), .A2(n19461), .B1(n20839), .B2(n20838), .O(
        n21361) );
  INV1S U23008 ( .I(n21361), .O(n20920) );
  XOR2HS U23009 ( .I1(n20840), .I2(n20920), .O(n20841) );
  XNR2HS U23010 ( .I1(n21200), .I2(n20841), .O(n20929) );
  INV1S U23011 ( .I(n20892), .O(n29451) );
  OR2 U23012 ( .I1(n23186), .I2(n20891), .O(n20844) );
  NR2 U23013 ( .I1(n13822), .I2(n23187), .O(n20842) );
  OAI112HS U23014 ( .C1(n29470), .C2(n23188), .A1(n20844), .B1(n20843), .O(
        n20846) );
  ND2S U23015 ( .I1(n29484), .I2(n20891), .O(n20845) );
  OAI112HS U23016 ( .C1(n29451), .C2(n21079), .A1(n20846), .B1(n20845), .O(
        n20848) );
  AOI22S U23017 ( .A1(n20899), .A2(n28533), .B1(n20848), .B2(n20847), .O(
        n20851) );
  OAI22S U23018 ( .A1(n23184), .A2(n20899), .B1(n22528), .B2(n21000), .O(
        n20850) );
  AOI22S U23019 ( .A1(n26015), .A2(n20903), .B1(n29505), .B2(n29519), .O(
        n20849) );
  OAI12HS U23020 ( .B1(n20851), .B2(n20850), .A1(n20849), .O(n20853) );
  INV1S U23021 ( .I(n20948), .O(n21007) );
  ND2S U23022 ( .I1(n21007), .I2(n22410), .O(n20852) );
  OAI112HS U23023 ( .C1(n23179), .C2(n29519), .A1(n20853), .B1(n20852), .O(
        n20854) );
  NR2 U23024 ( .I1(n22932), .I2(n20892), .O(n20862) );
  ND2S U23025 ( .I1(n29470), .I2(n13887), .O(n20856) );
  ND3S U23026 ( .I1(n20856), .I2(n22942), .I3(n22419), .O(n20860) );
  OAI22S U23027 ( .A1(n29489), .A2(n22416), .B1(n22415), .B2(n29448), .O(
        n20857) );
  AOI13HS U23028 ( .B1(n20860), .B2(n20859), .B3(n20858), .A1(n20857), .O(
        n20861) );
  OAI22S U23029 ( .A1(n20862), .A2(n20861), .B1(n22418), .B2(n21616), .O(
        n20865) );
  ND2S U23030 ( .I1(n20865), .I2(n20864), .O(n20868) );
  OA22 U23031 ( .A1(n19494), .A2(n22412), .B1(n22411), .B2(n29513), .O(n20867)
         );
  OAI22S U23032 ( .A1(n21254), .A2(n29519), .B1(n19461), .B2(n21259), .O(
        n20866) );
  AO12 U23033 ( .B1(n20868), .B2(n20867), .A1(n20866), .O(n20869) );
  OAI12HS U23034 ( .B1(n22410), .B2(n20855), .A1(n20869), .O(n21241) );
  OR2 U23035 ( .I1(n20991), .I2(n21241), .O(n20919) );
  INV1S U23036 ( .I(n20919), .O(n20871) );
  INV1S U23037 ( .I(n20991), .O(n21097) );
  INV1S U23038 ( .I(n21241), .O(n21292) );
  NR2 U23039 ( .I1(n21097), .I2(n21292), .O(n20870) );
  NR2 U23040 ( .I1(n20871), .I2(n20870), .O(n20914) );
  NR2 U23041 ( .I1(n22411), .I2(n17965), .O(n20885) );
  OAI22S U23042 ( .A1(n21403), .A2(n22415), .B1(n21407), .B2(n22418), .O(
        n20880) );
  ND2S U23043 ( .I1(n29491), .I2(n20891), .O(n20878) );
  ND2S U23044 ( .I1(n21394), .I2(n22417), .O(n20874) );
  ND3S U23045 ( .I1(n20874), .I2(n20873), .I3(n21643), .O(n20877) );
  OR2 U23046 ( .I1(n22417), .I2(n21394), .O(n20876) );
  OAI22S U23047 ( .A1(n22058), .A2(n20891), .B1(n20892), .B2(n22059), .O(
        n20875) );
  AOI13HS U23048 ( .B1(n20878), .B2(n20877), .B3(n20876), .A1(n20875), .O(
        n20879) );
  OAI22S U23049 ( .A1(n20880), .A2(n20879), .B1(n22062), .B2(n20899), .O(
        n20883) );
  OR2 U23050 ( .I1(n22412), .I2(n21412), .O(n20882) );
  OAI22S U23051 ( .A1(n22055), .A2(n20903), .B1(n29519), .B2(n22054), .O(
        n20881) );
  AOI12HS U23052 ( .B1(n20883), .B2(n20882), .A1(n20881), .O(n20884) );
  OAI22S U23053 ( .A1(n20885), .A2(n20884), .B1(n22053), .B2(n19461), .O(
        n20886) );
  OAI12HS U23054 ( .B1(n22410), .B2(n21449), .A1(n20886), .O(n21428) );
  NR2 U23055 ( .I1(n20891), .I2(n29497), .O(n20887) );
  NR2 U23056 ( .I1(n20895), .I2(n20887), .O(n20898) );
  NR2 U23057 ( .I1(n29470), .I2(n29475), .O(n20890) );
  AN2S U23058 ( .I1(n27893), .I2(n22419), .O(n20889) );
  ND2S U23059 ( .I1(n29475), .I2(n29470), .O(n20888) );
  OAI12HS U23060 ( .B1(n20890), .B2(n20889), .A1(n20888), .O(n20897) );
  ND2S U23061 ( .I1(n29497), .I2(n20891), .O(n20894) );
  ND2S U23062 ( .I1(n29455), .I2(n20892), .O(n20893) );
  OAI12HS U23063 ( .B1(n20895), .B2(n20894), .A1(n20893), .O(n20896) );
  AOI12HS U23064 ( .B1(n20898), .B2(n20897), .A1(n20896), .O(n20902) );
  NR2 U23065 ( .I1(n20899), .I2(n28527), .O(n20901) );
  ND2S U23066 ( .I1(n28527), .I2(n20899), .O(n20900) );
  OAI12H U23067 ( .B1(n20902), .B2(n20901), .A1(n20900), .O(n20906) );
  AN2 U23068 ( .I1(n19059), .I2(n20903), .O(n20904) );
  AOI12H U23069 ( .B1(n20906), .B2(n20905), .A1(n20904), .O(n20909) );
  NR2 U23070 ( .I1(n29519), .I2(n21416), .O(n20908) );
  ND2S U23071 ( .I1(n21416), .I2(n29519), .O(n20907) );
  OAI12H U23072 ( .B1(n20909), .B2(n20908), .A1(n20907), .O(n20912) );
  XNR2HS U23073 ( .I1(n21428), .I2(n21474), .O(n20913) );
  XNR2HS U23074 ( .I1(n20916), .I2(n20913), .O(n20928) );
  XNR2HS U23075 ( .I1(n20914), .I2(n20928), .O(n20915) );
  XNR2HS U23076 ( .I1(n20929), .I2(n20915), .O(n20935) );
  NR2 U23077 ( .I1(n21428), .I2(n21474), .O(n20917) );
  XNR2HS U23078 ( .I1(n20919), .I2(n20918), .O(n20923) );
  OR2 U23079 ( .I1(n20919), .I2(n20918), .O(n20927) );
  MAO222 U23080 ( .A1(n21128), .B1(n20921), .C1(n20920), .O(n20922) );
  MXL2HS U23081 ( .A(n20923), .B(n20927), .S(n20922), .OB(n20934) );
  INV1S U23082 ( .I(n20922), .O(n20925) );
  INV1S U23083 ( .I(n20923), .O(n20924) );
  NR2 U23084 ( .I1(n20925), .I2(n20924), .O(n20926) );
  AN3B2S U23085 ( .I1(n20927), .B1(n20926), .B2(n20934), .O(n20933) );
  INV1S U23086 ( .I(n20928), .O(n20931) );
  INV1S U23087 ( .I(n20929), .O(n20930) );
  ND2S U23088 ( .I1(n20931), .I2(n20930), .O(n20932) );
  OR2 U23089 ( .I1(n21386), .I2(n21388), .O(n21385) );
  NR2 U23090 ( .I1(n21641), .I2(n23187), .O(n20937) );
  NR2 U23091 ( .I1(n29467), .I2(n23188), .O(n20936) );
  OAI22S U23092 ( .A1(n13887), .A2(n21072), .B1(n20937), .B2(n20936), .O(
        n20939) );
  NR2 U23093 ( .I1(n21246), .I2(n21076), .O(n20938) );
  MOAI1S U23094 ( .A1(n20939), .A2(n20938), .B1(n21246), .B2(n23244), .O(
        n20940) );
  OAI12HS U23095 ( .B1(n21117), .B2(n21079), .A1(n20940), .O(n20941) );
  OAI12HS U23096 ( .B1(n20942), .B2(n13816), .A1(n20941), .O(n20943) );
  OAI12HS U23097 ( .B1(n21656), .B2(n21023), .A1(n20943), .O(n20946) );
  OA22 U23098 ( .A1(n23508), .A2(n21000), .B1(n23184), .B2(n21616), .O(n20945)
         );
  OAI22S U23099 ( .A1(n22920), .A2(n21088), .B1(n21081), .B2(n22922), .O(
        n20944) );
  AOI12HS U23100 ( .B1(n20946), .B2(n20945), .A1(n20944), .O(n20952) );
  OAI22S U23101 ( .A1(n20950), .A2(n20949), .B1(n20948), .B2(n20947), .O(
        n20951) );
  MOAI1 U23102 ( .A1(n20952), .A2(n20951), .B1(n23848), .B2(n20855), .O(n21285) );
  NR2 U23103 ( .I1(n28533), .I2(n24768), .O(n20954) );
  NR2 U23104 ( .I1(n28528), .I2(n26012), .O(n20955) );
  ND2P U23105 ( .I1(n21612), .I2(n21023), .O(n20956) );
  AOI12HS U23106 ( .B1(n20956), .B2(n26012), .A1(n24768), .O(n20953) );
  AOI22S U23107 ( .A1(n20954), .A2(n20955), .B1(n20953), .B2(n21081), .O(
        n20988) );
  INV1S U23108 ( .I(n20955), .O(n20959) );
  OAI112HS U23109 ( .C1(n28533), .C2(n20959), .A1(n20958), .B1(n24768), .O(
        n20960) );
  ND2 U23110 ( .I1(n20960), .I2(n21088), .O(n20987) );
  OAI22S U23111 ( .A1(n21596), .A2(n21081), .B1(n21612), .B2(n21023), .O(
        n20962) );
  NR2 U23112 ( .I1(n20962), .I2(n20961), .O(n20985) );
  NR2 U23113 ( .I1(n26638), .I2(n29462), .O(n20979) );
  AOI22S U23114 ( .A1(n21046), .A2(n13804), .B1(n20439), .B2(n21045), .O(
        n20967) );
  AOI22S U23115 ( .A1(n21063), .A2(n13835), .B1(n13847), .B2(n21059), .O(
        n20966) );
  AOI22S U23116 ( .A1(n21044), .A2(n13839), .B1(n13846), .B2(n21053), .O(
        n20965) );
  AOI22S U23117 ( .A1(n21049), .A2(n20963), .B1(n13791), .B2(n21038), .O(
        n20964) );
  AN4S U23118 ( .I1(n20967), .I2(n20966), .I3(n20965), .I4(n20964), .O(n20975)
         );
  AOI22S U23119 ( .A1(n21058), .A2(n20613), .B1(n17875), .B2(n21043), .O(
        n20973) );
  AOI22S U23120 ( .A1(n21054), .A2(n13830), .B1(n21062), .B2(n21040), .O(
        n20972) );
  AOI22S U23121 ( .A1(n21037), .A2(n20968), .B1(n17762), .B2(n21050), .O(
        n20971) );
  AOI22S U23122 ( .A1(n21060), .A2(n17928), .B1(n20969), .B2(n21039), .O(
        n20970) );
  AN4S U23123 ( .I1(n20973), .I2(n20972), .I3(n20971), .I4(n20970), .O(n20974)
         );
  ND2S U23124 ( .I1(n20975), .I2(n20974), .O(n20976) );
  MXL2HS U23125 ( .A(n22670), .B(n20977), .S(n13822), .OB(n27888) );
  ND2S U23126 ( .I1(n27891), .I2(n27888), .O(n20978) );
  MOAI1 U23127 ( .A1(n20979), .A2(n20978), .B1(n26638), .B2(n29462), .O(n20981) );
  ND2S U23128 ( .I1(n21079), .I2(n29444), .O(n20982) );
  ND2S U23129 ( .I1(n29485), .I2(n21076), .O(n20980) );
  ND3S U23130 ( .I1(n20981), .I2(n20982), .I3(n20980), .O(n20984) );
  ND3S U23131 ( .I1(n20982), .I2(n25391), .I3(n29484), .O(n20983) );
  ND3 U23132 ( .I1(n20988), .I2(n20987), .I3(n20986), .O(n20989) );
  ND2S U23133 ( .I1(n21394), .I2(n29462), .O(n20993) );
  ND3S U23134 ( .I1(n20993), .I2(n23427), .I3(n21643), .O(n20995) );
  OAI112HS U23135 ( .C1(n21399), .C2(n23186), .A1(n20995), .B1(n20994), .O(
        n20999) );
  ND2S U23136 ( .I1(n29443), .I2(n21403), .O(n20998) );
  ND2S U23137 ( .I1(n21399), .I2(n29484), .O(n20997) );
  OAI22S U23138 ( .A1(n21403), .A2(n23185), .B1(n21407), .B2(n23184), .O(
        n20996) );
  AOI13HS U23139 ( .B1(n20999), .B2(n20998), .B3(n20997), .A1(n20996), .O(
        n21003) );
  AN2S U23140 ( .I1(n21407), .I2(n28533), .O(n21002) );
  INV1S U23141 ( .I(n21000), .O(n21001) );
  ND2S U23142 ( .I1(n29505), .I2(n17965), .O(n21004) );
  ND3P U23143 ( .I1(n21005), .I2(n21004), .I3(n13935), .O(n21009) );
  AOI22S U23144 ( .A1(n21007), .A2(n22053), .B1(n21006), .B2(n22054), .O(
        n21008) );
  NR2 U23145 ( .I1(n21398), .I2(n21076), .O(n21010) );
  NR2 U23146 ( .I1(n29455), .I2(n21079), .O(n21016) );
  NR2 U23147 ( .I1(n21010), .I2(n21016), .O(n21019) );
  NR2 U23148 ( .I1(n29475), .I2(n21072), .O(n21013) );
  AN2S U23149 ( .I1(n27893), .I2(n27891), .O(n21012) );
  ND2 U23150 ( .I1(n21072), .I2(n29475), .O(n21011) );
  OAI12HS U23151 ( .B1(n21013), .B2(n21012), .A1(n21011), .O(n21018) );
  ND2S U23152 ( .I1(n21079), .I2(n29455), .O(n21014) );
  OAI12HS U23153 ( .B1(n21016), .B2(n21015), .A1(n21014), .O(n21017) );
  AOI12HS U23154 ( .B1(n21019), .B2(n21018), .A1(n21017), .O(n21035) );
  NR2P U23155 ( .I1(n23839), .I2(n21085), .O(n21029) );
  NR2 U23156 ( .I1(n21416), .I2(n21088), .O(n21020) );
  NR2P U23157 ( .I1(n21029), .I2(n21020), .O(n21032) );
  NR2 U23158 ( .I1(n21023), .I2(n28527), .O(n21021) );
  NR2 U23159 ( .I1(n21411), .I2(n21081), .O(n21026) );
  NR2 U23160 ( .I1(n21021), .I2(n21026), .O(n21022) );
  ND2P U23161 ( .I1(n21032), .I2(n21022), .O(n21034) );
  ND2S U23162 ( .I1(n28527), .I2(n21023), .O(n21025) );
  ND2S U23163 ( .I1(n21081), .I2(n21411), .O(n21024) );
  OAI12HS U23164 ( .B1(n21026), .B2(n21025), .A1(n21024), .O(n21031) );
  ND2S U23165 ( .I1(n21088), .I2(n21416), .O(n21028) );
  ND2S U23166 ( .I1(n21085), .I2(n23839), .O(n21027) );
  OAI12HS U23167 ( .B1(n21029), .B2(n21028), .A1(n21027), .O(n21030) );
  AOI12HS U23168 ( .B1(n21032), .B2(n21031), .A1(n21030), .O(n21033) );
  OAI12HP U23169 ( .B1(n21035), .B2(n21034), .A1(n21033), .O(n21477) );
  XOR2H U23170 ( .I1(n21425), .I2(n21477), .O(n21036) );
  XNR2H U23171 ( .I1(n21093), .I2(n21036), .O(n21092) );
  AOI22S U23172 ( .A1(n21038), .A2(n19914), .B1(n20263), .B2(n21037), .O(
        n21042) );
  AOI22S U23173 ( .A1(n21040), .A2(n13839), .B1(n13847), .B2(n21039), .O(
        n21041) );
  ND2S U23174 ( .I1(n21042), .I2(n21041), .O(n21069) );
  AOI22S U23175 ( .A1(n21044), .A2(n13846), .B1(n20187), .B2(n21043), .O(
        n21048) );
  AOI22S U23176 ( .A1(n21046), .A2(n20124), .B1(n17938), .B2(n21045), .O(
        n21047) );
  ND2S U23177 ( .I1(n21048), .I2(n21047), .O(n21068) );
  ND2S U23178 ( .I1(n21049), .I2(n17928), .O(n21052) );
  ND2S U23179 ( .I1(n21050), .I2(n13804), .O(n21051) );
  ND3S U23180 ( .I1(n21052), .I2(n21051), .I3(n13822), .O(n21057) );
  INV1S U23181 ( .I(n21053), .O(n21055) );
  MOAI1S U23182 ( .A1(n13844), .A2(n21055), .B1(n21054), .B2(n17762), .O(
        n21056) );
  NR2 U23183 ( .I1(n21057), .I2(n21056), .O(n21066) );
  AOI22S U23184 ( .A1(n21059), .A2(n13830), .B1(n17875), .B2(n21058), .O(
        n21065) );
  AOI22S U23185 ( .A1(n21063), .A2(n21062), .B1(n21061), .B2(n21060), .O(
        n21064) );
  ND3S U23186 ( .I1(n21066), .I2(n21065), .I3(n21064), .O(n21067) );
  NR3 U23187 ( .I1(n21069), .I2(n21068), .I3(n21067), .O(n21070) );
  NR2 U23188 ( .I1(n21329), .I2(n21070), .O(n21638) );
  INV1S U23189 ( .I(n26639), .O(n29464) );
  AOI22S U23190 ( .A1(n21071), .A2(n21638), .B1(n21072), .B2(n29464), .O(
        n21074) );
  NR2 U23191 ( .I1(n29464), .I2(n21072), .O(n21073) );
  MOAI1 U23192 ( .A1(n21074), .A2(n21073), .B1(n21076), .B2(n29486), .O(n21075) );
  OAI12HS U23193 ( .B1(n21076), .B2(n29486), .A1(n21075), .O(n21077) );
  OAI12HS U23194 ( .B1(n29445), .B2(n21079), .A1(n21078), .O(n21080) );
  NR2 U23195 ( .I1(n21597), .I2(n21081), .O(n21083) );
  AOI22S U23196 ( .A1(n21081), .A2(n21597), .B1(n21088), .B2(n29509), .O(
        n21082) );
  OAI12H U23197 ( .B1(n21084), .B2(n21083), .A1(n21082), .O(n21087) );
  OR2 U23198 ( .I1(n21460), .I2(n21085), .O(n21086) );
  OAI112H U23199 ( .C1(n29509), .C2(n21088), .A1(n21087), .B1(n21086), .O(
        n21089) );
  XNR2HS U23200 ( .I1(n21090), .I2(n21357), .O(n21103) );
  INV1S U23201 ( .I(n23841), .O(n21102) );
  ND2S U23202 ( .I1(n21477), .I2(n21425), .O(n21094) );
  ND2 U23203 ( .I1(n21094), .I2(n21093), .O(n21095) );
  OAI12HS U23204 ( .B1(n21477), .B2(n21425), .A1(n21095), .O(n21105) );
  NR2 U23205 ( .I1(n21096), .I2(n21357), .O(n23840) );
  INV1S U23206 ( .I(n21285), .O(n21098) );
  MAO222 U23207 ( .A1(n21199), .B1(n21098), .C1(n21097), .O(n21106) );
  ND3S U23208 ( .I1(n21105), .I2(n23840), .I3(n21106), .O(n21101) );
  XNR2HS U23209 ( .I1(n23840), .I2(n21105), .O(n21099) );
  INV1S U23210 ( .I(n21103), .O(n21111) );
  INV1S U23211 ( .I(n21104), .O(n21108) );
  NR2 U23212 ( .I1(n23840), .I2(n21105), .O(n21107) );
  OAI22S U23213 ( .A1(n21111), .A2(n21108), .B1(n21107), .B2(n21106), .O(
        n21112) );
  INV1S U23214 ( .I(n21109), .O(n21110) );
  MOAI1 U23215 ( .A1(n23841), .A2(n21112), .B1(n21111), .B2(n21110), .O(n21452) );
  OR2 U23216 ( .I1(n21641), .I2(n22670), .O(n21115) );
  INV1S U23217 ( .I(n29467), .O(n21113) );
  NR2 U23218 ( .I1(n21113), .I2(n26638), .O(n21114) );
  OAI22S U23219 ( .A1(n21115), .A2(n21114), .B1(n29467), .B2(n22668), .O(
        n21116) );
  OAI12HS U23220 ( .B1(n21246), .B2(n25391), .A1(n21116), .O(n21121) );
  OR2 U23221 ( .I1(n29448), .I2(n22671), .O(n21120) );
  OAI22S U23222 ( .A1(n21117), .A2(n27262), .B1(n28528), .B2(n21656), .O(
        n21118) );
  AOI13HS U23223 ( .B1(n21121), .B2(n21120), .B3(n21119), .A1(n21118), .O(
        n21124) );
  OAI22S U23224 ( .A1(n19494), .A2(n22663), .B1(n22669), .B2(n21616), .O(
        n21123) );
  OAI12HS U23225 ( .B1(n21124), .B2(n21123), .A1(n21122), .O(n21126) );
  OAI112HS U23226 ( .C1(n22662), .C2(n29513), .A1(n21126), .B1(n21125), .O(
        n21127) );
  OAI12HS U23227 ( .B1(n21237), .B2(n23845), .A1(n21127), .O(n21291) );
  MAO222 U23228 ( .A1(n21199), .B1(n21291), .C1(n21128), .O(n21155) );
  NR2 U23229 ( .I1(n29445), .I2(n27262), .O(n21135) );
  NR2 U23230 ( .I1(n29486), .I2(n25391), .O(n21129) );
  NR2 U23231 ( .I1(n21135), .I2(n21129), .O(n21138) );
  NR2 U23232 ( .I1(n29464), .I2(n26638), .O(n21132) );
  INV1S U23233 ( .I(n21638), .O(n27889) );
  INV1S U23234 ( .I(n27888), .O(n21637) );
  ND2S U23235 ( .I1(n26638), .I2(n29464), .O(n21130) );
  OAI12HS U23236 ( .B1(n21132), .B2(n21131), .A1(n21130), .O(n21137) );
  ND2S U23237 ( .I1(n25391), .I2(n29486), .O(n21134) );
  ND2S U23238 ( .I1(n27262), .I2(n29445), .O(n21133) );
  OAI12HS U23239 ( .B1(n21135), .B2(n21134), .A1(n21133), .O(n21136) );
  AOI12HS U23240 ( .B1(n21138), .B2(n21137), .A1(n21136), .O(n21153) );
  NR2 U23241 ( .I1(n21460), .I2(n23845), .O(n21146) );
  NR2 U23242 ( .I1(n29509), .I2(n24768), .O(n21139) );
  NR2 U23243 ( .I1(n21146), .I2(n21139), .O(n21150) );
  NR2 U23244 ( .I1(n21613), .I2(n28528), .O(n21140) );
  NR2 U23245 ( .I1(n21597), .I2(n26012), .O(n21144) );
  NR2 U23246 ( .I1(n21140), .I2(n21144), .O(n21141) );
  ND2S U23247 ( .I1(n21150), .I2(n21141), .O(n21152) );
  ND2S U23248 ( .I1(n28528), .I2(n21613), .O(n21143) );
  ND2S U23249 ( .I1(n26012), .I2(n21597), .O(n21142) );
  OAI12HS U23250 ( .B1(n21144), .B2(n21143), .A1(n21142), .O(n21149) );
  ND2S U23251 ( .I1(n24768), .I2(n29509), .O(n21147) );
  ND2S U23252 ( .I1(n23845), .I2(n21460), .O(n21145) );
  OAI12HS U23253 ( .B1(n21147), .B2(n21146), .A1(n21145), .O(n21148) );
  AOI12HS U23254 ( .B1(n21150), .B2(n21149), .A1(n21148), .O(n21151) );
  OAI12H U23255 ( .B1(n21153), .B2(n21152), .A1(n21151), .O(n21360) );
  OR2 U23256 ( .I1(n21154), .I2(n21360), .O(n21202) );
  INV1S U23257 ( .I(n21202), .O(n23843) );
  ND2S U23258 ( .I1(n21155), .I2(n23843), .O(n21210) );
  INV1S U23259 ( .I(n21210), .O(n21198) );
  INV1S U23260 ( .I(n21155), .O(n21156) );
  INV1S U23261 ( .I(n21212), .O(n21197) );
  ND2S U23262 ( .I1(n27893), .I2(n21637), .O(n21157) );
  MAO222 U23263 ( .A1(n21157), .B1(n26638), .C1(n29475), .O(n21158) );
  NR2 U23264 ( .I1(n28528), .I2(n28527), .O(n21162) );
  NR2 U23265 ( .I1(n29455), .I2(n27262), .O(n21159) );
  NR2 U23266 ( .I1(n21162), .I2(n21159), .O(n21164) );
  ND2 U23267 ( .I1(n28527), .I2(n28528), .O(n21160) );
  OAI12HS U23268 ( .B1(n21162), .B2(n21161), .A1(n21160), .O(n21163) );
  AOI12HS U23269 ( .B1(n21165), .B2(n21164), .A1(n21163), .O(n21176) );
  NR2 U23270 ( .I1(n21411), .I2(n26012), .O(n21166) );
  NR2 U23271 ( .I1(n21416), .I2(n24768), .O(n21170) );
  NR2 U23272 ( .I1(n21166), .I2(n21170), .O(n21167) );
  OR2 U23273 ( .I1(n23839), .I2(n23845), .O(n21172) );
  ND2S U23274 ( .I1(n21167), .I2(n21172), .O(n21175) );
  ND2 U23275 ( .I1(n26012), .I2(n21411), .O(n21169) );
  OAI12HS U23276 ( .B1(n21170), .B2(n21169), .A1(n21168), .O(n21173) );
  AOI12HS U23277 ( .B1(n21173), .B2(n21172), .A1(n21171), .O(n21174) );
  OAI12H U23278 ( .B1(n21176), .B2(n21175), .A1(n21174), .O(n21471) );
  NR2 U23279 ( .I1(n21194), .I2(n21471), .O(n21196) );
  NR2 U23280 ( .I1(n22670), .I2(n21177), .O(n21178) );
  NR2 U23281 ( .I1(n22730), .I2(n21178), .O(n21180) );
  INV1S U23282 ( .I(n21394), .O(n29469) );
  AOI12HS U23283 ( .B1(n21178), .B2(n26638), .A1(n29469), .O(n21179) );
  OAI22S U23284 ( .A1(n21180), .A2(n21179), .B1(n22667), .B2(n21399), .O(
        n21183) );
  AOI22S U23285 ( .A1(n21399), .A2(n29485), .B1(n21403), .B2(n29444), .O(
        n21182) );
  OR2 U23286 ( .I1(n22663), .I2(n21412), .O(n21184) );
  OAI12HS U23287 ( .B1(n21403), .B2(n22671), .A1(n21184), .O(n21181) );
  AOI12HS U23288 ( .B1(n21183), .B2(n21182), .A1(n21181), .O(n21188) );
  ND2S U23289 ( .I1(n21407), .I2(n21612), .O(n21186) );
  INV1S U23290 ( .I(n21184), .O(n21185) );
  NR2 U23291 ( .I1(n21186), .I2(n21185), .O(n21187) );
  MOAI1 U23292 ( .A1(n21188), .A2(n21187), .B1(n28528), .B2(n21618), .O(n21190) );
  ND2S U23293 ( .I1(n29508), .I2(n17965), .O(n21189) );
  OAI112HS U23294 ( .C1(n26012), .C2(n21601), .A1(n21190), .B1(n21189), .O(
        n21193) );
  AOI22H U23295 ( .A1(n21457), .A2(n21449), .B1(n21193), .B2(n21192), .O(
        n21438) );
  INV1S U23296 ( .I(n21438), .O(n21195) );
  MOAI1 U23297 ( .A1(n21196), .A2(n21195), .B1(n21471), .B2(n21194), .O(n21211) );
  MXL2HS U23298 ( .A(n21198), .B(n21197), .S(n21211), .OB(n21209) );
  XNR2HS U23299 ( .I1(n21291), .I2(n21199), .O(n21201) );
  INV1S U23300 ( .I(n21360), .O(n21204) );
  OAI12HS U23301 ( .B1(n21204), .B2(n21203), .A1(n21202), .O(n21214) );
  XOR2HS U23302 ( .I1(n21438), .I2(n21471), .O(n21205) );
  XNR2HS U23303 ( .I1(n21206), .I2(n21205), .O(n21216) );
  ND2S U23304 ( .I1(n21211), .I2(n21210), .O(n21213) );
  OAI12H U23305 ( .B1(n21216), .B2(n21215), .A1(n21214), .O(n23844) );
  AO12T U23306 ( .B1(n21453), .B2(n21452), .A1(n21456), .O(n21458) );
  XOR2HS U23307 ( .I1(n21220), .I2(n21285), .O(n21244) );
  INV2 U23308 ( .I(n29486), .O(n25392) );
  OR2 U23309 ( .I1(n21641), .I2(n21221), .O(n21223) );
  NR2 U23310 ( .I1(n13887), .I2(n26639), .O(n21222) );
  OAI22S U23311 ( .A1(n21223), .A2(n21222), .B1(n29467), .B2(n21333), .O(
        n21224) );
  OAI12HS U23312 ( .B1(n21246), .B2(n25392), .A1(n21224), .O(n21227) );
  ND2S U23313 ( .I1(n21330), .I2(n21225), .O(n21226) );
  OAI112HS U23314 ( .C1(n21228), .C2(n29448), .A1(n21227), .B1(n21226), .O(
        n21230) );
  ND2S U23315 ( .I1(n29445), .I2(n29448), .O(n21229) );
  AOI22S U23316 ( .A1(n21656), .A2(n21231), .B1(n21230), .B2(n21229), .O(
        n21233) );
  NR2 U23317 ( .I1(n21656), .I2(n28531), .O(n21232) );
  MOAI1 U23318 ( .A1(n21233), .A2(n21232), .B1(n21340), .B2(n21245), .O(n21235) );
  ND2S U23319 ( .I1(n29509), .I2(n29513), .O(n21234) );
  OAI112HS U23320 ( .C1(n22922), .C2(n26013), .A1(n21235), .B1(n21234), .O(
        n21240) );
  AOI22S U23321 ( .A1(n21238), .A2(n21237), .B1(n21345), .B2(n21254), .O(
        n21239) );
  AOI22S U23322 ( .A1(n21460), .A2(n20855), .B1(n21240), .B2(n21239), .O(
        n21304) );
  XNR2HS U23323 ( .I1(n21304), .I2(n21241), .O(n21242) );
  XNR2HS U23324 ( .I1(n21291), .I2(n21242), .O(n21293) );
  INV1S U23325 ( .I(n21293), .O(n21243) );
  XNR2HS U23326 ( .I1(n21244), .I2(n21243), .O(n21282) );
  OAI22S U23327 ( .A1(n29513), .A2(n22054), .B1(n22055), .B2(n19494), .O(
        n21256) );
  OR2 U23328 ( .I1(n21245), .I2(n21412), .O(n21250) );
  ND3S U23329 ( .I1(n21250), .I2(n21656), .I3(n21407), .O(n21253) );
  OAI22S U23330 ( .A1(n29489), .A2(n22058), .B1(n22061), .B2(n29467), .O(
        n21248) );
  MAOI1 U23331 ( .A1(n22942), .A2(n21643), .B1(n13887), .B2(n21394), .O(n21247) );
  OAI22S U23332 ( .A1(n21248), .A2(n21247), .B1(n21246), .B2(n21399), .O(
        n21249) );
  OAI12HS U23333 ( .B1(n22059), .B2(n29448), .A1(n21249), .O(n21251) );
  AOI22S U23334 ( .A1(n21618), .A2(n21616), .B1(n21253), .B2(n21252), .O(
        n21255) );
  OAI22S U23335 ( .A1(n21256), .A2(n21255), .B1(n21254), .B2(n17965), .O(
        n21257) );
  OAI12HS U23336 ( .B1(n21449), .B2(n21259), .A1(n21258), .O(n21424) );
  INV1S U23337 ( .I(n21424), .O(n21426) );
  ND2S U23338 ( .I1(n27893), .I2(n21260), .O(n21261) );
  MAO222 U23339 ( .A1(n21261), .B1(n29467), .C1(n29475), .O(n21262) );
  MAO222 U23340 ( .A1(n21262), .B1(n29489), .C1(n29497), .O(n21269) );
  NR2 U23341 ( .I1(n29448), .I2(n29455), .O(n21263) );
  NR2 U23342 ( .I1(n21616), .I2(n28527), .O(n21266) );
  NR2 U23343 ( .I1(n21263), .I2(n21266), .O(n21268) );
  ND2S U23344 ( .I1(n29455), .I2(n29448), .O(n21265) );
  ND2S U23345 ( .I1(n28527), .I2(n21616), .O(n21264) );
  OAI12HS U23346 ( .B1(n21266), .B2(n21265), .A1(n21264), .O(n21267) );
  AOI12HS U23347 ( .B1(n21269), .B2(n21268), .A1(n21267), .O(n21276) );
  OR2S U23348 ( .I1(n19494), .I2(n19059), .O(n21270) );
  OR2 U23349 ( .I1(n29513), .I2(n21416), .O(n21273) );
  ND2S U23350 ( .I1(n21270), .I2(n21273), .O(n21275) );
  AN2S U23351 ( .I1(n19059), .I2(n19494), .O(n21272) );
  AOI12HS U23352 ( .B1(n21273), .B2(n21272), .A1(n21271), .O(n21274) );
  OAI12HS U23353 ( .B1(n21276), .B2(n21275), .A1(n21274), .O(n21279) );
  OR2 U23354 ( .I1(n20855), .I2(n23839), .O(n21278) );
  AO12T U23355 ( .B1(n21279), .B2(n21278), .A1(n21277), .O(n21478) );
  XOR2HS U23356 ( .I1(n21280), .I2(n21478), .O(n21281) );
  XNR2HS U23357 ( .I1(n21426), .I2(n21281), .O(n21294) );
  XNR2HS U23358 ( .I1(n21282), .I2(n21294), .O(n21303) );
  NR2 U23359 ( .I1(n21424), .I2(n21478), .O(n21284) );
  MOAI1 U23360 ( .A1(n21284), .A2(n21283), .B1(n21478), .B2(n21424), .O(n21287) );
  INV1S U23361 ( .I(n21287), .O(n21290) );
  OR2 U23362 ( .I1(n21286), .I2(n21285), .O(n21288) );
  INV1S U23363 ( .I(n21288), .O(n21289) );
  OAI12HS U23364 ( .B1(n21290), .B2(n21289), .A1(n21298), .O(n21299) );
  INV1S U23365 ( .I(n21304), .O(n21359) );
  MAO222 U23366 ( .A1(n21292), .B1(n21359), .C1(n21291), .O(n21297) );
  ND2S U23367 ( .I1(n21294), .I2(n21293), .O(n21296) );
  ND2S U23368 ( .I1(n21296), .I2(n21298), .O(n21295) );
  AOI12HS U23369 ( .B1(n21299), .B2(n21297), .A1(n21295), .O(n21302) );
  INV1S U23370 ( .I(n21296), .O(n21301) );
  MXL2HS U23371 ( .A(n21299), .B(n21298), .S(n21297), .OB(n21300) );
  XOR2HS U23372 ( .I1(n21304), .I2(n21360), .O(n21305) );
  XNR2HS U23373 ( .I1(n21361), .I2(n21305), .O(n21351) );
  NR2 U23374 ( .I1(n27263), .I2(n29455), .O(n21312) );
  NR2 U23375 ( .I1(n25392), .I2(n29497), .O(n21306) );
  NR2 U23376 ( .I1(n21312), .I2(n21306), .O(n21315) );
  NR2 U23377 ( .I1(n26639), .I2(n29475), .O(n21309) );
  ND2S U23378 ( .I1(n29475), .I2(n26639), .O(n21308) );
  OAI12HS U23379 ( .B1(n21309), .B2(n21307), .A1(n21308), .O(n21314) );
  ND2S U23380 ( .I1(n29497), .I2(n25392), .O(n21311) );
  ND2S U23381 ( .I1(n29455), .I2(n27263), .O(n21310) );
  OAI12HS U23382 ( .B1(n21312), .B2(n21311), .A1(n21310), .O(n21313) );
  AOI12HS U23383 ( .B1(n21315), .B2(n21314), .A1(n21313), .O(n21325) );
  NR2 U23384 ( .I1(n26013), .I2(n19059), .O(n21320) );
  NR2 U23385 ( .I1(n28531), .I2(n28527), .O(n21316) );
  NR2 U23386 ( .I1(n21320), .I2(n21316), .O(n21317) );
  INV1S U23387 ( .I(n29509), .O(n24769) );
  ND2S U23388 ( .I1(n21317), .I2(n13923), .O(n21324) );
  ND2S U23389 ( .I1(n28527), .I2(n28531), .O(n21319) );
  ND2S U23390 ( .I1(n19059), .I2(n26013), .O(n21318) );
  OAI12HS U23391 ( .B1(n21320), .B2(n21319), .A1(n21318), .O(n21322) );
  AOI12HS U23392 ( .B1(n21322), .B2(n13923), .A1(n21321), .O(n21323) );
  OAI12HS U23393 ( .B1(n21325), .B2(n21324), .A1(n21323), .O(n21328) );
  OR2 U23394 ( .I1(n23846), .I2(n23839), .O(n21327) );
  AO12T U23395 ( .B1(n21328), .B2(n21327), .A1(n21326), .O(n21476) );
  MOAI1 U23396 ( .A1(n29491), .A2(n25392), .B1(n21403), .B2(n29445), .O(n21338) );
  NR2 U23397 ( .I1(n26639), .I2(n22061), .O(n21332) );
  ND2S U23398 ( .I1(n22060), .I2(n21329), .O(n21331) );
  MOAI1S U23399 ( .A1(n21332), .A2(n21331), .B1(n21330), .B2(n22058), .O(
        n21335) );
  NR2 U23400 ( .I1(n21333), .I2(n21394), .O(n21334) );
  NR2 U23401 ( .I1(n21335), .I2(n21334), .O(n21337) );
  INV1 U23402 ( .I(n21403), .O(n29450) );
  MOAI1 U23403 ( .A1(n21338), .A2(n21337), .B1(n29450), .B2(n21336), .O(n21339) );
  AOI22S U23404 ( .A1(n21412), .A2(n21597), .B1(n17965), .B2(n29509), .O(
        n21343) );
  AOI22S U23405 ( .A1(n22053), .A2(n21346), .B1(n21345), .B2(n22054), .O(
        n21347) );
  AOI22HP U23406 ( .A1(n21449), .A2(n21460), .B1(n21348), .B2(n21347), .O(
        n21436) );
  XNR2HS U23407 ( .I1(n21350), .I2(n21357), .O(n21368) );
  ND2S U23408 ( .I1(n21352), .I2(n21351), .O(n21366) );
  OAI12H U23409 ( .B1(n21369), .B2(n21368), .A1(n21366), .O(n21380) );
  NR2 U23410 ( .I1(n21353), .I2(n21476), .O(n21355) );
  INV1S U23411 ( .I(n21436), .O(n21354) );
  MOAI1 U23412 ( .A1(n21355), .A2(n21354), .B1(n21476), .B2(n21353), .O(n21374) );
  ND2S U23413 ( .I1(n21374), .I2(n21377), .O(n21358) );
  ND2S U23414 ( .I1(n21380), .I2(n21358), .O(n21365) );
  INV3CK U23415 ( .I(n21377), .O(n21363) );
  NR2 U23416 ( .I1(n21359), .I2(n21360), .O(n21362) );
  XNR2HS U23417 ( .I1(n21364), .I2(n21374), .O(n21367) );
  ND2S U23418 ( .I1(n21365), .I2(n21367), .O(n21383) );
  NR2 U23419 ( .I1(n21367), .I2(n21366), .O(n21373) );
  INV1S U23420 ( .I(n21368), .O(n21371) );
  INV1S U23421 ( .I(n21369), .O(n21370) );
  XNR2HS U23422 ( .I1(n21371), .I2(n21370), .O(n21372) );
  NR2 U23423 ( .I1(n21373), .I2(n21372), .O(n21382) );
  INV1S U23424 ( .I(n21375), .O(n21376) );
  NR2 U23425 ( .I1(n21377), .I2(n21376), .O(n21378) );
  OR2T U23426 ( .I1(n21381), .I2(n21380), .O(n28530) );
  ND3P U23427 ( .I1(n21383), .I2(n21382), .I3(n28530), .O(n21459) );
  ND3HT U23428 ( .I1(n21450), .I2(n21384), .I3(n21459), .O(n21387) );
  NR2F U23429 ( .I1(n21385), .I2(n21387), .O(n29516) );
  ND2F U23430 ( .I1(n21446), .I2(n29516), .O(n29504) );
  INV1 U23431 ( .I(n21386), .O(n21389) );
  NR2T U23432 ( .I1(n21389), .I2(n21387), .O(n29502) );
  INV1S U23433 ( .I(n21387), .O(n21390) );
  AN2T U23434 ( .I1(n21390), .I2(n13934), .O(n29521) );
  AOI22S U23435 ( .A1(n21392), .A2(n29502), .B1(n29521), .B2(n21391), .O(
        n21466) );
  INV2 U23436 ( .I(n21393), .O(n21430) );
  AN2S U23437 ( .I1(n27893), .I2(n21643), .O(n21397) );
  NR2 U23438 ( .I1(n21394), .I2(n29475), .O(n21396) );
  ND2S U23439 ( .I1(n29475), .I2(n21394), .O(n21395) );
  OAI12HS U23440 ( .B1(n21397), .B2(n21396), .A1(n21395), .O(n21402) );
  AN2S U23441 ( .I1(n29497), .I2(n21399), .O(n21400) );
  NR2 U23442 ( .I1(n29455), .I2(n21403), .O(n21405) );
  ND2S U23443 ( .I1(n21403), .I2(n29455), .O(n21404) );
  OAI12H U23444 ( .B1(n21406), .B2(n21405), .A1(n21404), .O(n21410) );
  AN2 U23445 ( .I1(n28527), .I2(n21407), .O(n21408) );
  AOI12H U23446 ( .B1(n21410), .B2(n21409), .A1(n21408), .O(n21415) );
  NR2 U23447 ( .I1(n21412), .I2(n21411), .O(n21414) );
  OAI12H U23448 ( .B1(n21415), .B2(n21414), .A1(n21413), .O(n21419) );
  OR2 U23449 ( .I1(n21416), .I2(n17965), .O(n21418) );
  NR2 U23450 ( .I1(n21449), .I2(n23839), .O(n21421) );
  XOR2HS U23451 ( .I1(n21428), .I2(n21470), .O(n21423) );
  XNR2HS U23452 ( .I1(n21430), .I2(n21423), .O(n21445) );
  XNR2HS U23453 ( .I1(n21425), .I2(n21424), .O(n21434) );
  ND2S U23454 ( .I1(n21445), .I2(n21434), .O(n21439) );
  INV1S U23455 ( .I(n21425), .O(n21427) );
  NR2 U23456 ( .I1(n21427), .I2(n21426), .O(n21432) );
  MOAI1S U23457 ( .A1(n21470), .A2(n21430), .B1(n21429), .B2(n21428), .O(
        n21431) );
  ND2S U23458 ( .I1(n21431), .I2(n21432), .O(n21444) );
  OAI12HS U23459 ( .B1(n21432), .B2(n21431), .A1(n21444), .O(n21441) );
  XNR3 U23460 ( .I1(n21433), .I2(n21439), .I3(n21441), .O(n21448) );
  OAI12HS U23461 ( .B1(n21445), .B2(n21434), .A1(n21439), .O(n21437) );
  XOR4S U23462 ( .I1(n21438), .I2(n21437), .I3(n21436), .I4(n21435), .O(n21443) );
  INV1S U23463 ( .I(n21439), .O(n21440) );
  ND3S U23464 ( .I1(n21441), .I2(n21440), .I3(n21444), .O(n21442) );
  OAI112HS U23465 ( .C1(n21445), .C2(n21444), .A1(n21443), .B1(n21442), .O(
        n21447) );
  NR3HT U23466 ( .I1(n21448), .I2(n21447), .I3(n21446), .O(n29518) );
  INV1S U23467 ( .I(n21449), .O(n21464) );
  ND3P U23468 ( .I1(n21451), .I2(n21450), .I3(n21459), .O(n29514) );
  INV1S U23469 ( .I(n21453), .O(n21454) );
  NR3HP U23470 ( .I1(n21456), .I2(n21455), .I3(n21454), .O(n29506) );
  AOI22S U23471 ( .A1(n29507), .A2(n21457), .B1(n29506), .B2(n23848), .O(
        n21462) );
  NR2P U23472 ( .I1(n21459), .I2(n21458), .O(n29510) );
  ND2S U23473 ( .I1(n29510), .I2(n21460), .O(n21461) );
  OAI112HS U23474 ( .C1(n29514), .C2(n20855), .A1(n21462), .B1(n21461), .O(
        n21463) );
  AOI13HS U23475 ( .B1(n29518), .B2(n21464), .B3(n29516), .A1(n21463), .O(
        n21465) );
  NR2 U23476 ( .I1(n21471), .I2(n21472), .O(n21469) );
  INV1S U23477 ( .I(n21470), .O(n21468) );
  MOAI1 U23478 ( .A1(n21469), .A2(n21468), .B1(n21471), .B2(n21472), .O(n21496) );
  XOR2HS U23479 ( .I1(n21481), .I2(n21496), .O(n21488) );
  XOR2HS U23480 ( .I1(n21477), .I2(n21474), .O(n21475) );
  XNR2HS U23481 ( .I1(n21478), .I2(n21475), .O(n21489) );
  OAI12HS U23482 ( .B1(n13909), .B2(n21476), .A1(n21481), .O(n21490) );
  OAI12HS U23483 ( .B1(n21492), .B2(n21489), .A1(n21490), .O(n21482) );
  NR2 U23484 ( .I1(n21477), .I2(n21478), .O(n21480) );
  MOAI1S U23485 ( .A1(n21480), .A2(n21479), .B1(n21478), .B2(n21477), .O(
        n21483) );
  ND2S U23486 ( .I1(n21482), .I2(n21483), .O(n21495) );
  INV1S U23487 ( .I(n21481), .O(n21497) );
  INV1S U23488 ( .I(n21482), .O(n21485) );
  INV1S U23489 ( .I(n21483), .O(n21484) );
  OAI112HS U23490 ( .C1(n21496), .C2(n21497), .A1(n21485), .B1(n21484), .O(
        n21486) );
  ND2 U23491 ( .I1(n21495), .I2(n21486), .O(n21487) );
  XNR2HS U23492 ( .I1(n21488), .I2(n21487), .O(n21500) );
  INV1S U23493 ( .I(n21489), .O(n21491) );
  XNR2HS U23494 ( .I1(n21491), .I2(n21490), .O(n21494) );
  INV1S U23495 ( .I(n21492), .O(n21493) );
  XNR2HS U23496 ( .I1(n21494), .I2(n21493), .O(n21499) );
  INV1S U23497 ( .I(n21495), .O(n21498) );
  ND3S U23498 ( .I1(n21500), .I2(n21499), .I3(n28536), .O(n21502) );
  AN2 U23499 ( .I1(n21502), .I2(n23770), .O(n29527) );
  INV1S U23500 ( .I(A67_shift[7]), .O(n21505) );
  INV1S U23501 ( .I(n23839), .O(n21504) );
  NR2P U23502 ( .I1(n29526), .I2(n21502), .O(n29525) );
  INV1S U23503 ( .I(n29525), .O(n21503) );
  OAI222S U23504 ( .A1(n13907), .A2(n21651), .B1(n23770), .B2(n21505), .C1(
        n21504), .C2(n21503), .O(n11485) );
  NR2 U23505 ( .I1(n21513), .I2(n21514), .O(n21565) );
  NR2 U23506 ( .I1(n21584), .I2(n21565), .O(n21516) );
  NR2 U23507 ( .I1(n21509), .I2(n21510), .O(n23433) );
  NR2 U23508 ( .I1(rgb_value[0]), .I2(rgb_value[16]), .O(n23459) );
  INV1S U23509 ( .I(rgb_value[8]), .O(n21506) );
  ND2S U23510 ( .I1(rgb_value[16]), .I2(rgb_value[0]), .O(n23460) );
  OAI12HS U23511 ( .B1(n23459), .B2(n21506), .A1(n23460), .O(n23453) );
  ND2S U23512 ( .I1(n21507), .I2(rgb_value[9]), .O(n23451) );
  INV1S U23513 ( .I(n23451), .O(n21508) );
  AOI12HS U23514 ( .B1(n13928), .B2(n23453), .A1(n21508), .O(n23437) );
  ND2S U23515 ( .I1(n21510), .I2(n21509), .O(n23434) );
  OAI12HS U23516 ( .B1(n23433), .B2(n23437), .A1(n23434), .O(n21568) );
  ND2S U23517 ( .I1(n21512), .I2(n21511), .O(n21585) );
  ND2S U23518 ( .I1(n21514), .I2(n21513), .O(n21566) );
  OAI12HS U23519 ( .B1(n21565), .B2(n21585), .A1(n21566), .O(n21515) );
  AOI12HS U23520 ( .B1(n21516), .B2(n21568), .A1(n21515), .O(n21531) );
  NR2 U23521 ( .I1(n21519), .I2(n21520), .O(n21537) );
  NR2 U23522 ( .I1(n21537), .I2(n21540), .O(n21533) );
  ND2S U23523 ( .I1(n21533), .I2(n13930), .O(n21525) );
  ND2S U23524 ( .I1(n21518), .I2(n21517), .O(n21556) );
  ND2S U23525 ( .I1(n21520), .I2(n21519), .O(n21538) );
  OAI12HS U23526 ( .B1(n21537), .B2(n21556), .A1(n21538), .O(n21532) );
  ND2S U23527 ( .I1(n21522), .I2(n21521), .O(n21530) );
  INV1S U23528 ( .I(n21530), .O(n21523) );
  AOI12HS U23529 ( .B1(n21532), .B2(n13930), .A1(n21523), .O(n21524) );
  OAI12HS U23530 ( .B1(n21531), .B2(n21525), .A1(n21524), .O(n21526) );
  INV1S U23531 ( .I(n21528), .O(n21529) );
  ND2S U23532 ( .I1(n13930), .I2(n21530), .O(n21535) );
  INV1S U23533 ( .I(n21531), .O(n21558) );
  AOI12HS U23534 ( .B1(n21558), .B2(n21533), .A1(n21532), .O(n21534) );
  XOR2HS U23535 ( .I1(n21535), .I2(n21534), .O(n21551) );
  INV1 U23536 ( .I(n21551), .O(n21550) );
  NR2 U23537 ( .I1(n21529), .I2(n21550), .O(n21536) );
  INV1S U23538 ( .I(n21537), .O(n21539) );
  ND2S U23539 ( .I1(n21539), .I2(n21538), .O(n21543) );
  INV1S U23540 ( .I(n21540), .O(n21557) );
  INV1S U23541 ( .I(n21556), .O(n21541) );
  AOI12HS U23542 ( .B1(n21558), .B2(n21557), .A1(n21541), .O(n21542) );
  XOR2HS U23543 ( .I1(n21543), .I2(n21542), .O(n21561) );
  NR2 U23544 ( .I1(n21560), .I2(n21550), .O(n21544) );
  NR2 U23545 ( .I1(n21544), .I2(n21528), .O(n21548) );
  INV1S U23546 ( .I(n21545), .O(n21546) );
  INV1S U23547 ( .I(gray_avg[7]), .O(n21549) );
  AOI22S U23548 ( .A1(gray_avg[7]), .A2(n21550), .B1(n21549), .B2(n21551), .O(
        n21555) );
  XOR2HS U23549 ( .I1(n21560), .I2(n21551), .O(n21552) );
  INV1S U23550 ( .I(n21552), .O(n21553) );
  MXL2HS U23551 ( .A(n21553), .B(n21552), .S(gray_avg[7]), .OB(n21554) );
  MXL2HS U23552 ( .A(n21555), .B(n21554), .S(gray_avg[6]), .OB(n21573) );
  ND2S U23553 ( .I1(n21557), .I2(n21556), .O(n21559) );
  XNR2HS U23554 ( .I1(n21559), .I2(n21558), .O(n21579) );
  INV1S U23555 ( .I(n21579), .O(n21578) );
  INV1 U23556 ( .I(gray_avg[6]), .O(n21562) );
  MOAI1 U23557 ( .A1(n21561), .A2(n21562), .B1(n21562), .B2(n21561), .O(n21571) );
  NR2 U23558 ( .I1(n21578), .I2(n21563), .O(n21564) );
  INV1S U23559 ( .I(n21565), .O(n21567) );
  ND2S U23560 ( .I1(n21567), .I2(n21566), .O(n21570) );
  INV1S U23561 ( .I(n21568), .O(n21587) );
  OAI12HS U23562 ( .B1(n21587), .B2(n21584), .A1(n21585), .O(n21569) );
  XNR2HS U23563 ( .I1(n21570), .I2(n21569), .O(n21590) );
  INV1S U23564 ( .I(n21590), .O(n21589) );
  NR2 U23565 ( .I1(n21589), .I2(n21578), .O(n21572) );
  NR2 U23566 ( .I1(n21572), .I2(n21571), .O(n21576) );
  INV1S U23567 ( .I(n21573), .O(n21574) );
  INV1S U23568 ( .I(gray_avg[5]), .O(n21577) );
  AOI22S U23569 ( .A1(gray_avg[5]), .A2(n21578), .B1(n21577), .B2(n21579), .O(
        n21583) );
  AN2B1S U23570 ( .I1(n21578), .B1(n21589), .O(n21581) );
  XOR2HS U23571 ( .I1(n21589), .I2(n21579), .O(n21580) );
  MXL2HS U23572 ( .A(n21581), .B(n21580), .S(gray_avg[5]), .OB(n21582) );
  MXL2HS U23573 ( .A(n21583), .B(n21582), .S(gray_avg[4]), .OB(n23440) );
  INV1S U23574 ( .I(n21584), .O(n21586) );
  ND2S U23575 ( .I1(n21586), .I2(n21585), .O(n21588) );
  XOR2HS U23576 ( .I1(n21588), .I2(n21587), .O(n23446) );
  INV1S U23577 ( .I(n23446), .O(n23445) );
  INV1 U23578 ( .I(gray_avg[4]), .O(n21591) );
  INV1S U23579 ( .I(n23438), .O(n21592) );
  NR2 U23580 ( .I1(n23445), .I2(n21592), .O(n21593) );
  MOAI1 U23581 ( .A1(n29504), .A2(n21595), .B1(n29502), .B2(n21594), .O(n21605) );
  AOI22S U23582 ( .A1(n29507), .A2(n21596), .B1(n29506), .B2(n26015), .O(
        n21599) );
  ND2S U23583 ( .I1(n29510), .I2(n21597), .O(n21598) );
  OAI112HS U23584 ( .C1(n29514), .C2(n19494), .A1(n21599), .B1(n21598), .O(
        n21600) );
  AOI13HS U23585 ( .B1(n29518), .B2(n21601), .B3(n29516), .A1(n21600), .O(
        n21604) );
  OR3B2 U23586 ( .I1(n21605), .B1(n21604), .B2(n21603), .O(n21606) );
  INV1S U23587 ( .I(n21606), .O(n21609) );
  INV1S U23588 ( .I(A67_shift[5]), .O(n21608) );
  INV1S U23589 ( .I(n19059), .O(n21607) );
  MOAI1 U23590 ( .A1(n29504), .A2(n21611), .B1(n29502), .B2(n21610), .O(n21622) );
  AOI22S U23591 ( .A1(n29507), .A2(n21612), .B1(n29506), .B2(n28533), .O(
        n21615) );
  ND2S U23592 ( .I1(n29510), .I2(n21613), .O(n21614) );
  OAI112HS U23593 ( .C1(n29514), .C2(n21616), .A1(n21615), .B1(n21614), .O(
        n21617) );
  AOI13HS U23594 ( .B1(n29518), .B2(n21618), .B3(n29516), .A1(n21617), .O(
        n21621) );
  OR3B2 U23595 ( .I1(n21622), .B1(n21621), .B2(n21620), .O(n21623) );
  INV1S U23596 ( .I(n21623), .O(n21626) );
  INV1S U23597 ( .I(A67_shift[4]), .O(n21625) );
  INV1S U23598 ( .I(n28527), .O(n21624) );
  XNR2HS U23599 ( .I1(n21628), .I2(n21627), .O(n21629) );
  XNR2HS U23600 ( .I1(n21630), .I2(n21629), .O(PE_N71) );
  XOR2HS U23601 ( .I1(n21632), .I2(n21631), .O(n21633) );
  XNR2HS U23602 ( .I1(n21634), .I2(n21633), .O(PE_N58) );
  INV1S U23603 ( .I(n29504), .O(n21636) );
  ND2S U23604 ( .I1(n21636), .I2(n21635), .O(n21647) );
  AOI22S U23605 ( .A1(n29507), .A2(n21637), .B1(n29506), .B2(n27891), .O(
        n21640) );
  ND2S U23606 ( .I1(n29510), .I2(n21638), .O(n21639) );
  OAI112HS U23607 ( .C1(n29514), .C2(n21641), .A1(n21640), .B1(n21639), .O(
        n21642) );
  AOI13HS U23608 ( .B1(n29518), .B2(n21643), .B3(n29516), .A1(n21642), .O(
        n21646) );
  AOI22S U23609 ( .A1(n21644), .A2(n29502), .B1(n29521), .B2(n22419), .O(
        n21645) );
  ND3 U23610 ( .I1(n21647), .I2(n21646), .I3(n21645), .O(n21648) );
  INV1S U23611 ( .I(n21648), .O(n21652) );
  INV1S U23612 ( .I(n29527), .O(n21651) );
  INV1S U23613 ( .I(A67_shift[0]), .O(n21650) );
  INV1S U23614 ( .I(template_store[24]), .O(n22397) );
  INV1S U23615 ( .I(n21653), .O(n22302) );
  NR2 U23616 ( .I1(n22397), .I2(n22302), .O(n21668) );
  INV1S U23617 ( .I(template_store[27]), .O(n22323) );
  NR2 U23618 ( .I1(n22323), .I2(n13815), .O(n21667) );
  INV1S U23619 ( .I(template_store[26]), .O(n21714) );
  NR2 U23620 ( .I1(n21714), .I2(n13765), .O(n21671) );
  INV1S U23621 ( .I(template_store[30]), .O(n22348) );
  NR2 U23622 ( .I1(n22348), .I2(n20735), .O(n21670) );
  INV1S U23623 ( .I(template_store[29]), .O(n22333) );
  NR2 U23624 ( .I1(n22333), .I2(n22331), .O(n21674) );
  INV1S U23625 ( .I(template_store[28]), .O(n21713) );
  NR2 U23626 ( .I1(n21713), .I2(n13813), .O(n21673) );
  INV1S U23627 ( .I(template_store[25]), .O(n22325) );
  NR2 U23628 ( .I1(n22325), .I2(n13765), .O(n21662) );
  NR2 U23629 ( .I1(n22333), .I2(n20735), .O(n21661) );
  NR2 U23630 ( .I1(n22325), .I2(n22322), .O(n21665) );
  NR2 U23631 ( .I1(n22397), .I2(n22322), .O(n21682) );
  NR2 U23632 ( .I1(n22323), .I2(n13813), .O(n21681) );
  NR2 U23633 ( .I1(n22397), .I2(n13765), .O(n21676) );
  NR2 U23634 ( .I1(n21713), .I2(n20735), .O(n21675) );
  NR2 U23635 ( .I1(n21713), .I2(n22331), .O(n21679) );
  NR2 U23636 ( .I1(n21714), .I2(n13815), .O(n21678) );
  HA1 U23637 ( .A(n21662), .B(n21661), .C(n21672), .S(n21677) );
  NR2 U23638 ( .I1(n22325), .I2(n22302), .O(n22354) );
  NR2 U23639 ( .I1(n21713), .I2(n13815), .O(n22353) );
  NR2 U23640 ( .I1(n22323), .I2(n13765), .O(n22327) );
  INV1S U23641 ( .I(template_store[31]), .O(n22332) );
  NR2 U23642 ( .I1(n22332), .I2(n20735), .O(n22326) );
  FA1 U23643 ( .A(n21665), .B(n21664), .CI(n21663), .CO(n22374), .S(n21683) );
  NR2 U23644 ( .I1(n22348), .I2(n22331), .O(n22351) );
  NR2 U23645 ( .I1(n22397), .I2(n22324), .O(n22350) );
  HA1 U23646 ( .A(n21671), .B(n21670), .C(n22349), .S(n21666) );
  NR2 U23647 ( .I1(n21714), .I2(n22322), .O(n22341) );
  NR2 U23648 ( .I1(n22333), .I2(n13813), .O(n22340) );
  FA1 U23649 ( .A(n21674), .B(n21673), .CI(n21672), .CO(n22339), .S(n21684) );
  NR2 U23650 ( .I1(n22323), .I2(n22331), .O(n21688) );
  NR2 U23651 ( .I1(n22325), .I2(n13815), .O(n21687) );
  HA1 U23652 ( .A(n21676), .B(n21675), .C(n21680), .S(n21686) );
  FA1 U23653 ( .A(n21679), .B(n21678), .CI(n21677), .CO(n21663), .S(n21700) );
  FA1 U23654 ( .A(n21685), .B(n21684), .CI(n21683), .CO(n22378), .S(n22380) );
  FA1 U23655 ( .A(n21688), .B(n21687), .CI(n21686), .CO(n21701), .S(n22384) );
  NR2 U23656 ( .I1(n21714), .I2(n13813), .O(n21698) );
  NR2 U23657 ( .I1(n22323), .I2(n20735), .O(n21690) );
  NR2 U23658 ( .I1(n21714), .I2(n22331), .O(n21689) );
  NR2 U23659 ( .I1(n22325), .I2(n13813), .O(n21695) );
  NR2 U23660 ( .I1(n22397), .I2(n13815), .O(n21694) );
  NR2 U23661 ( .I1(n21714), .I2(n20735), .O(n21692) );
  NR2 U23662 ( .I1(n22325), .I2(n22331), .O(n21691) );
  NR2 U23663 ( .I1(n22397), .I2(n13813), .O(n22390) );
  NR2 U23664 ( .I1(n22325), .I2(n20735), .O(n22409) );
  NR2 U23665 ( .I1(n22397), .I2(n22331), .O(n22408) );
  HA1 U23666 ( .A(n21692), .B(n21691), .C(n21693), .S(n22388) );
  FA1 U23667 ( .A(n21701), .B(n21700), .CI(n21699), .CO(n22381), .S(n21719) );
  NR2 U23668 ( .I1(n21720), .I2(n21719), .O(n21702) );
  MOAI1 U23669 ( .A1(n21703), .A2(n21702), .B1(n21719), .B2(n21720), .O(n22379) );
  NR2 U23670 ( .I1(n22332), .I2(n13765), .O(n21706) );
  NR2 U23671 ( .I1(n22333), .I2(n22302), .O(n21705) );
  NR2 U23672 ( .I1(n21713), .I2(n22324), .O(n21704) );
  NR2 U23673 ( .I1(n22348), .I2(n22302), .O(n22305) );
  NR2 U23674 ( .I1(n22332), .I2(n22322), .O(n22304) );
  NR2 U23675 ( .I1(n22333), .I2(n22324), .O(n22303) );
  NR2 U23676 ( .I1(n22348), .I2(n22322), .O(n21709) );
  NR2 U23677 ( .I1(n22348), .I2(n13765), .O(n21712) );
  NR2 U23678 ( .I1(n21713), .I2(n22302), .O(n21711) );
  NR2 U23679 ( .I1(n22332), .I2(n13815), .O(n21710) );
  FA1S U23680 ( .A(n21706), .B(n21705), .CI(n21704), .CO(n22311), .S(n21707)
         );
  NR2 U23681 ( .I1(n22333), .I2(n22322), .O(n21717) );
  NR2 U23682 ( .I1(n22323), .I2(n22324), .O(n21716) );
  NR2 U23683 ( .I1(n22333), .I2(n13765), .O(n22330) );
  NR2 U23684 ( .I1(n22323), .I2(n22302), .O(n22329) );
  NR2 U23685 ( .I1(n22348), .I2(n13815), .O(n22328) );
  FA1S U23686 ( .A(n21709), .B(n21708), .CI(n21707), .CO(n22309), .S(n22406)
         );
  FA1S U23687 ( .A(n21712), .B(n21711), .CI(n21710), .CO(n21708), .S(n22360)
         );
  NR2 U23688 ( .I1(n21713), .I2(n22322), .O(n22344) );
  NR2 U23689 ( .I1(n21714), .I2(n22324), .O(n22343) );
  NR2 U23690 ( .I1(n21713), .I2(n13765), .O(n22335) );
  NR2 U23691 ( .I1(n21714), .I2(n22302), .O(n22334) );
  FA1S U23692 ( .A(n21717), .B(n21716), .CI(n21715), .CO(n22407), .S(n22358)
         );
  XOR2HS U23693 ( .I1(n22312), .I2(n22313), .O(n21718) );
  XNR2HS U23694 ( .I1(n21718), .I2(n22315), .O(PE_N92) );
  XNR2HS U23695 ( .I1(n21720), .I2(n21719), .O(n21721) );
  XNR2HS U23696 ( .I1(n21722), .I2(n21721), .O(PE_N85) );
  FA1 U23697 ( .A(n21725), .B(n21724), .CI(n21723), .CO(n23556), .S(PE_N67) );
  NR2 U23698 ( .I1(n21727), .I2(n21238), .O(n21757) );
  NR2 U23699 ( .I1(n21730), .I2(n21238), .O(n21733) );
  NR2 U23700 ( .I1(n21727), .I2(n21729), .O(n21732) );
  NR2 U23701 ( .I1(n21727), .I2(n21726), .O(n21739) );
  NR2 U23702 ( .I1(n21728), .I2(n21238), .O(n21738) );
  NR2 U23703 ( .I1(n21730), .I2(n21729), .O(n21737) );
  FA1S U23704 ( .A(n21733), .B(n21732), .CI(n21731), .CO(n21756), .S(n21760)
         );
  FA1S U23705 ( .A(n21736), .B(n21735), .CI(n21734), .CO(n21745), .S(n21740)
         );
  FA1S U23706 ( .A(n21739), .B(n21738), .CI(n21737), .CO(n21731), .S(n21744)
         );
  FA1S U23707 ( .A(n21742), .B(n21741), .CI(n21740), .CO(n21743), .S(n21747)
         );
  FA1S U23708 ( .A(n21745), .B(n21744), .CI(n21743), .CO(n21759), .S(n21763)
         );
  FA1S U23709 ( .A(n21748), .B(n21747), .CI(n21746), .CO(n21762), .S(n21750)
         );
  INV1S U23710 ( .I(n21750), .O(n21754) );
  INV1S U23711 ( .I(n21751), .O(n21753) );
  FA1 U23712 ( .A(n21757), .B(n21756), .CI(n21755), .CO(PE_N63), .S(PE_N62) );
  FA1 U23713 ( .A(n21760), .B(n21759), .CI(n21758), .CO(n21755), .S(PE_N61) );
  FA1 U23714 ( .A(n21763), .B(n21762), .CI(n21761), .CO(n21758), .S(PE_N60) );
  FA1 U23715 ( .A(n21766), .B(n21765), .CI(n21764), .CO(n15907), .S(n21798) );
  FA1 U23716 ( .A(n21772), .B(n21771), .CI(n21770), .CO(n21794), .S(n21796) );
  ND2S U23717 ( .I1(n21802), .I2(n21801), .O(mult_x_431_n10) );
  NR2 U23718 ( .I1(n21801), .I2(n21802), .O(mult_x_431_n9) );
  FA1 U23719 ( .A(n21778), .B(n21777), .CI(n21776), .CO(mult_x_431_n11), .S(
        PE_N55) );
  FA1 U23720 ( .A(n21781), .B(n21780), .CI(n21779), .CO(n21776), .S(PE_N54) );
  FA1 U23721 ( .A(n21784), .B(n21783), .CI(n21782), .CO(n15920), .S(PE_N52) );
  FA1 U23722 ( .A(n21787), .B(n21786), .CI(n21785), .CO(n21782), .S(PE_N51) );
  FA1 U23723 ( .A(n21795), .B(n21794), .CI(n21793), .CO(n21632), .S(
        mult_x_431_n39) );
  FA1 U23724 ( .A(n21798), .B(n21797), .CI(n21796), .CO(mult_x_431_n48), .S(
        n21802) );
  NR2 U23725 ( .I1(n21800), .I2(n21799), .O(PE_N48) );
  INV1S U23726 ( .I(template_store[15]), .O(n21915) );
  NR2 U23727 ( .I1(n21915), .I2(n13812), .O(n21806) );
  INV1S U23728 ( .I(template_store[14]), .O(n21920) );
  NR2 U23729 ( .I1(n21920), .I2(n13812), .O(n21947) );
  NR2 U23730 ( .I1(n21915), .I2(n21918), .O(n21946) );
  INV1S U23731 ( .I(template_store[13]), .O(n21919) );
  NR2 U23732 ( .I1(n21919), .I2(n13812), .O(n21953) );
  NR2 U23733 ( .I1(n21920), .I2(n21918), .O(n21952) );
  NR2 U23734 ( .I1(n21915), .I2(n13814), .O(n21951) );
  OR2S U23735 ( .I1(n21806), .I2(n21807), .O(n22051) );
  ND2S U23736 ( .I1(n21807), .I2(n21806), .O(n22049) );
  ND2S U23737 ( .I1(n22051), .I2(n22049), .O(n21975) );
  INV1S U23738 ( .I(template_store[11]), .O(n21916) );
  NR2 U23739 ( .I1(n21916), .I2(n21914), .O(n21828) );
  INV1S U23740 ( .I(template_store[9]), .O(n21872) );
  NR2 U23741 ( .I1(n21872), .I2(n21918), .O(n21827) );
  INV2 U23742 ( .I(n21809), .O(n22043) );
  NR2 U23743 ( .I1(n21915), .I2(n22043), .O(n21825) );
  INV1S U23744 ( .I(template_store[8]), .O(n22044) );
  NR2 U23745 ( .I1(n22044), .I2(n13812), .O(n21824) );
  NR2 U23746 ( .I1(n22044), .I2(n21918), .O(n21883) );
  INV1S U23747 ( .I(template_store[12]), .O(n21917) );
  NR2 U23748 ( .I1(n21917), .I2(n21871), .O(n21855) );
  INV1S U23749 ( .I(template_store[10]), .O(n21850) );
  NR2 U23750 ( .I1(n21850), .I2(n21910), .O(n21854) );
  NR2 U23751 ( .I1(n21917), .I2(n22043), .O(n21857) );
  NR2 U23752 ( .I1(n21850), .I2(n21849), .O(n21856) );
  NR2 U23753 ( .I1(n21850), .I2(n21914), .O(n21817) );
  NR2 U23754 ( .I1(n21872), .I2(n13814), .O(n21816) );
  NR2 U23755 ( .I1(n21920), .I2(n22043), .O(n21814) );
  NR2 U23756 ( .I1(n21917), .I2(n21849), .O(n21813) );
  NR2 U23757 ( .I1(n21919), .I2(n21849), .O(n21820) );
  NR2 U23758 ( .I1(n21850), .I2(n13814), .O(n21819) );
  HA1 U23759 ( .A(n21814), .B(n21813), .C(n21818), .S(n21815) );
  FA1S U23760 ( .A(n21817), .B(n21816), .CI(n21815), .CO(n21822), .S(n21881)
         );
  NR2 U23761 ( .I1(n21920), .I2(n21871), .O(n21831) );
  NR2 U23762 ( .I1(n21917), .I2(n21910), .O(n21830) );
  NR2 U23763 ( .I1(n21919), .I2(n21871), .O(n21886) );
  NR2 U23764 ( .I1(n21916), .I2(n21910), .O(n21885) );
  NR2 U23765 ( .I1(n21919), .I2(n22043), .O(n21852) );
  NR2 U23766 ( .I1(n21916), .I2(n21849), .O(n21851) );
  NR2 U23767 ( .I1(n21850), .I2(n21918), .O(n21848) );
  FA1S U23768 ( .A(n21820), .B(n21819), .CI(n21818), .CO(n21847), .S(n21823)
         );
  NR2 U23769 ( .I1(n21917), .I2(n21914), .O(n21845) );
  NR2 U23770 ( .I1(n21916), .I2(n13814), .O(n21844) );
  NR2 U23771 ( .I1(n21920), .I2(n21849), .O(n21839) );
  NR2 U23772 ( .I1(n21872), .I2(n13812), .O(n21838) );
  FA1S U23773 ( .A(n21823), .B(n21822), .CI(n21821), .CO(n21833), .S(n21899)
         );
  NR2 U23774 ( .I1(n21915), .I2(n21871), .O(n21837) );
  NR2 U23775 ( .I1(n21919), .I2(n21910), .O(n21836) );
  FA1S U23776 ( .A(n21828), .B(n21827), .CI(n21826), .CO(n21841), .S(n21901)
         );
  FA1S U23777 ( .A(n21831), .B(n21830), .CI(n21829), .CO(n21840), .S(n21821)
         );
  NR2 U23778 ( .I1(n21904), .I2(n21905), .O(n22009) );
  FA1S U23779 ( .A(n21834), .B(n21833), .CI(n21832), .CO(n21906), .S(n21905)
         );
  NR2 U23780 ( .I1(n21919), .I2(n21914), .O(n21932) );
  FA1S U23781 ( .A(n21837), .B(n21836), .CI(n21835), .CO(n21931), .S(n21842)
         );
  NR2 U23782 ( .I1(n21915), .I2(n21849), .O(n21923) );
  NR2 U23783 ( .I1(n21917), .I2(n13814), .O(n21922) );
  FA1S U23784 ( .A(n21842), .B(n21841), .CI(n21840), .CO(n21940), .S(n21832)
         );
  NR2 U23785 ( .I1(n21850), .I2(n13812), .O(n21913) );
  NR2 U23786 ( .I1(n21916), .I2(n21918), .O(n21912) );
  NR2 U23787 ( .I1(n21920), .I2(n21910), .O(n21911) );
  FA1S U23788 ( .A(n21845), .B(n21844), .CI(n21843), .CO(n21937), .S(n21846)
         );
  FA1S U23789 ( .A(n21848), .B(n21847), .CI(n21846), .CO(n21936), .S(n21834)
         );
  NR2 U23790 ( .I1(n21906), .I2(n21907), .O(n22003) );
  NR2 U23791 ( .I1(n22009), .I2(n22003), .O(n21909) );
  NR2 U23792 ( .I1(n21916), .I2(n21871), .O(n21863) );
  NR2 U23793 ( .I1(n21916), .I2(n22043), .O(n21865) );
  NR2 U23794 ( .I1(n21872), .I2(n21849), .O(n21864) );
  NR2 U23795 ( .I1(n21850), .I2(n21871), .O(n21868) );
  NR2 U23796 ( .I1(n22044), .I2(n21910), .O(n21867) );
  NR2 U23797 ( .I1(n22044), .I2(n21849), .O(n21870) );
  NR2 U23798 ( .I1(n21850), .I2(n22043), .O(n21869) );
  NR2 U23799 ( .I1(n21872), .I2(n21914), .O(n21889) );
  NR2 U23800 ( .I1(n22044), .I2(n13814), .O(n21888) );
  HA1 U23801 ( .A(n21852), .B(n21851), .C(n21884), .S(n21887) );
  FA1S U23802 ( .A(n21855), .B(n21854), .CI(n21853), .CO(n21882), .S(n21891)
         );
  NR2 U23803 ( .I1(n22044), .I2(n21914), .O(n21860) );
  NR2 U23804 ( .I1(n21872), .I2(n21910), .O(n21859) );
  HA1 U23805 ( .A(n21857), .B(n21856), .C(n21853), .S(n21858) );
  NR2 U23806 ( .I1(n21879), .I2(n21880), .O(n22023) );
  FA1S U23807 ( .A(n21860), .B(n21859), .CI(n21858), .CO(n21890), .S(n21876)
         );
  FA1S U23808 ( .A(n21863), .B(n21862), .CI(n21861), .CO(n21879), .S(n21877)
         );
  OR2 U23809 ( .I1(n21876), .I2(n21877), .O(n22029) );
  FA1S U23810 ( .A(n21868), .B(n21867), .CI(n21866), .CO(n21861), .S(n21875)
         );
  NR2 U23811 ( .I1(n21874), .I2(n21875), .O(n22032) );
  NR2 U23812 ( .I1(n22044), .I2(n21871), .O(n22045) );
  NR2 U23813 ( .I1(n21872), .I2(n22043), .O(n22046) );
  ND2S U23814 ( .I1(n22045), .I2(n22046), .O(n22047) );
  INV1S U23815 ( .I(n22047), .O(n22042) );
  NR2 U23816 ( .I1(n21872), .I2(n21871), .O(n22038) );
  ND2S U23817 ( .I1(n22037), .I2(n22038), .O(n22039) );
  INV1S U23818 ( .I(n22039), .O(n21873) );
  NR2 U23819 ( .I1(n22042), .I2(n21873), .O(n22036) );
  ND2S U23820 ( .I1(n21875), .I2(n21874), .O(n22033) );
  OAI12HS U23821 ( .B1(n22032), .B2(n22036), .A1(n22033), .O(n22031) );
  INV1S U23822 ( .I(n22028), .O(n21878) );
  AOI12HS U23823 ( .B1(n22029), .B2(n22031), .A1(n21878), .O(n22027) );
  OAI12HS U23824 ( .B1(n22023), .B2(n22027), .A1(n22024), .O(n22021) );
  FA1S U23825 ( .A(n21883), .B(n21882), .CI(n21881), .CO(n21900), .S(n21893)
         );
  FA1S U23826 ( .A(n21886), .B(n21885), .CI(n21884), .CO(n21829), .S(n21898)
         );
  FA1S U23827 ( .A(n21889), .B(n21888), .CI(n21887), .CO(n21897), .S(n21892)
         );
  FA1S U23828 ( .A(n21892), .B(n21891), .CI(n21890), .CO(n21896), .S(n21880)
         );
  OR2 U23829 ( .I1(n21893), .I2(n21894), .O(n22020) );
  INV1S U23830 ( .I(n22019), .O(n21895) );
  AOI12HS U23831 ( .B1(n22021), .B2(n22020), .A1(n21895), .O(n22018) );
  FA1S U23832 ( .A(n21898), .B(n21897), .CI(n21896), .CO(n21902), .S(n21894)
         );
  FA1S U23833 ( .A(n21901), .B(n21900), .CI(n21899), .CO(n21904), .S(n21903)
         );
  NR2 U23834 ( .I1(n21902), .I2(n21903), .O(n22014) );
  OAI12HS U23835 ( .B1(n22018), .B2(n22014), .A1(n22015), .O(n22006) );
  OAI12HS U23836 ( .B1(n22003), .B2(n22010), .A1(n22004), .O(n21908) );
  NR2 U23837 ( .I1(n21920), .I2(n21914), .O(n21929) );
  NR2 U23838 ( .I1(n21915), .I2(n21910), .O(n21928) );
  FA1S U23839 ( .A(n21913), .B(n21912), .CI(n21911), .CO(n21927), .S(n21938)
         );
  NR2 U23840 ( .I1(n21915), .I2(n21914), .O(n21956) );
  NR2 U23841 ( .I1(n21916), .I2(n13812), .O(n21926) );
  NR2 U23842 ( .I1(n21917), .I2(n21918), .O(n21925) );
  NR2 U23843 ( .I1(n21919), .I2(n13814), .O(n21924) );
  NR2 U23844 ( .I1(n21917), .I2(n13812), .O(n21950) );
  NR2 U23845 ( .I1(n21919), .I2(n21918), .O(n21949) );
  NR2 U23846 ( .I1(n21920), .I2(n13814), .O(n21948) );
  FA1S U23847 ( .A(n21923), .B(n21922), .CI(n21921), .CO(n21935), .S(n21930)
         );
  FA1S U23848 ( .A(n21926), .B(n21925), .CI(n21924), .CO(n21955), .S(n21934)
         );
  FA1S U23849 ( .A(n21929), .B(n21928), .CI(n21927), .CO(n21962), .S(n21933)
         );
  FA1S U23850 ( .A(n21932), .B(n21931), .CI(n21930), .CO(n21944), .S(n21941)
         );
  FA1S U23851 ( .A(n21935), .B(n21934), .CI(n21933), .CO(n21960), .S(n21943)
         );
  FA1S U23852 ( .A(n21938), .B(n21937), .CI(n21936), .CO(n21942), .S(n21939)
         );
  NR2 U23853 ( .I1(n21965), .I2(n21966), .O(n21991) );
  FA1S U23854 ( .A(n21944), .B(n21943), .CI(n21942), .CO(n21966), .S(n21964)
         );
  NR2 U23855 ( .I1(n21963), .I2(n21964), .O(n21995) );
  NR2 U23856 ( .I1(n21991), .I2(n21995), .O(n21979) );
  FA1S U23857 ( .A(n21947), .B(n21946), .CI(n21945), .CO(n21807), .S(n21969)
         );
  FA1S U23858 ( .A(n21950), .B(n21949), .CI(n21948), .CO(n21959), .S(n21954)
         );
  FA1S U23859 ( .A(n21953), .B(n21952), .CI(n21951), .CO(n21945), .S(n21958)
         );
  FA1S U23860 ( .A(n21956), .B(n21955), .CI(n21954), .CO(n21957), .S(n21961)
         );
  NR2 U23861 ( .I1(n21969), .I2(n21970), .O(n21976) );
  FA1S U23862 ( .A(n21959), .B(n21958), .CI(n21957), .CO(n21970), .S(n21967)
         );
  FA1S U23863 ( .A(n21962), .B(n21961), .CI(n21960), .CO(n21968), .S(n21965)
         );
  NR2 U23864 ( .I1(n21967), .I2(n21968), .O(n21983) );
  NR2 U23865 ( .I1(n21976), .I2(n21983), .O(n21972) );
  ND2 U23866 ( .I1(n21966), .I2(n21965), .O(n21992) );
  OAI12HS U23867 ( .B1(n21991), .B2(n21999), .A1(n21992), .O(n21980) );
  ND2 U23868 ( .I1(n21968), .I2(n21967), .O(n21987) );
  OAI12HS U23869 ( .B1(n21987), .B2(n21976), .A1(n21977), .O(n21971) );
  AOI12HS U23870 ( .B1(n21980), .B2(n21972), .A1(n21971), .O(n21973) );
  OAI12HS U23871 ( .B1(n21994), .B2(n21974), .A1(n21973), .O(n22052) );
  XNR2HS U23872 ( .I1(n21975), .I2(n22052), .O(PE_N126) );
  INV1S U23873 ( .I(n21976), .O(n21978) );
  ND2S U23874 ( .I1(n21978), .I2(n21977), .O(n21986) );
  INV1S U23875 ( .I(n21979), .O(n21982) );
  INV1S U23876 ( .I(n21980), .O(n21981) );
  OAI12HS U23877 ( .B1(n21994), .B2(n21982), .A1(n21981), .O(n21989) );
  INV1S U23878 ( .I(n21983), .O(n21988) );
  INV1S U23879 ( .I(n21987), .O(n21984) );
  XOR2HS U23880 ( .I1(n21986), .I2(n21985), .O(PE_N125) );
  ND2S U23881 ( .I1(n21988), .I2(n21987), .O(n21990) );
  XNR2HS U23882 ( .I1(n21990), .I2(n21989), .O(PE_N124) );
  INV1S U23883 ( .I(n21991), .O(n21993) );
  INV1S U23884 ( .I(n21995), .O(n22000) );
  INV1S U23885 ( .I(n21999), .O(n21996) );
  AOI12HS U23886 ( .B1(n22001), .B2(n22000), .A1(n21996), .O(n21997) );
  XOR2HS U23887 ( .I1(n21998), .I2(n21997), .O(PE_N123) );
  XNR2HS U23888 ( .I1(n22002), .I2(n22001), .O(PE_N122) );
  INV1S U23889 ( .I(n22003), .O(n22005) );
  INV1S U23890 ( .I(n22006), .O(n22013) );
  OAI12HS U23891 ( .B1(n22013), .B2(n22009), .A1(n22010), .O(n22007) );
  XNR2HS U23892 ( .I1(n22008), .I2(n22007), .O(PE_N121) );
  INV1S U23893 ( .I(n22009), .O(n22011) );
  ND2S U23894 ( .I1(n22011), .I2(n22010), .O(n22012) );
  XOR2HS U23895 ( .I1(n22013), .I2(n22012), .O(PE_N120) );
  INV1S U23896 ( .I(n22014), .O(n22016) );
  ND2S U23897 ( .I1(n22016), .I2(n22015), .O(n22017) );
  XOR2HS U23898 ( .I1(n22018), .I2(n22017), .O(PE_N119) );
  ND2S U23899 ( .I1(n22020), .I2(n22019), .O(n22022) );
  XNR2HS U23900 ( .I1(n22022), .I2(n22021), .O(PE_N118) );
  INV1S U23901 ( .I(n22023), .O(n22025) );
  ND2S U23902 ( .I1(n22025), .I2(n22024), .O(n22026) );
  XOR2HS U23903 ( .I1(n22027), .I2(n22026), .O(PE_N117) );
  ND2S U23904 ( .I1(n22029), .I2(n22028), .O(n22030) );
  XNR2HS U23905 ( .I1(n22031), .I2(n22030), .O(PE_N116) );
  INV1S U23906 ( .I(n22032), .O(n22034) );
  ND2S U23907 ( .I1(n22034), .I2(n22033), .O(n22035) );
  XOR2HS U23908 ( .I1(n22036), .I2(n22035), .O(PE_N115) );
  OR2S U23909 ( .I1(n22038), .I2(n22037), .O(n22040) );
  ND2S U23910 ( .I1(n22040), .I2(n22039), .O(n22041) );
  XNR2HS U23911 ( .I1(n22042), .I2(n22041), .O(PE_N114) );
  NR2 U23912 ( .I1(n22044), .I2(n22043), .O(PE_N112) );
  OR2S U23913 ( .I1(n22046), .I2(n22045), .O(n22048) );
  AN2S U23914 ( .I1(n22048), .I2(n22047), .O(PE_N113) );
  INV1S U23915 ( .I(n22049), .O(n22050) );
  AO12 U23916 ( .B1(n22052), .B2(n22051), .A1(n22050), .O(PE_N127) );
  INV1S U23917 ( .I(template_store[7]), .O(n22166) );
  NR2 U23918 ( .I1(n22166), .I2(n13809), .O(n22056) );
  INV1S U23919 ( .I(template_store[6]), .O(n22169) );
  NR2 U23920 ( .I1(n22169), .I2(n13809), .O(n22199) );
  NR2 U23921 ( .I1(n22166), .I2(n22171), .O(n22198) );
  NR2 U23922 ( .I1(n22166), .I2(n22168), .O(n22205) );
  INV1S U23923 ( .I(template_store[5]), .O(n22172) );
  NR2 U23924 ( .I1(n22172), .I2(n13809), .O(n22204) );
  NR2 U23925 ( .I1(n22169), .I2(n22171), .O(n22203) );
  OR2S U23926 ( .I1(n22056), .I2(n22057), .O(n22300) );
  ND2S U23927 ( .I1(n22057), .I2(n22056), .O(n22298) );
  ND2S U23928 ( .I1(n22300), .I2(n22298), .O(n22227) );
  INV1S U23929 ( .I(template_store[4]), .O(n22170) );
  NR2 U23930 ( .I1(n22170), .I2(n22118), .O(n22065) );
  INV1S U23931 ( .I(template_store[3]), .O(n22167) );
  NR2 U23932 ( .I1(n22167), .I2(n22162), .O(n22064) );
  NR2 U23933 ( .I1(n22169), .I2(n17195), .O(n22067) );
  NR2 U23934 ( .I1(n22172), .I2(n22121), .O(n22066) );
  INV1S U23935 ( .I(template_store[0]), .O(n22293) );
  NR2 U23936 ( .I1(n22293), .I2(n22171), .O(n22135) );
  NR2 U23937 ( .I1(n22293), .I2(n22168), .O(n22106) );
  INV1S U23938 ( .I(template_store[1]), .O(n22122) );
  NR2 U23939 ( .I1(n22122), .I2(n13810), .O(n22105) );
  NR2 U23940 ( .I1(n22170), .I2(n17195), .O(n22103) );
  NR2 U23941 ( .I1(n22167), .I2(n22121), .O(n22102) );
  FA1S U23942 ( .A(n22065), .B(n22064), .CI(n22063), .CO(n22153), .S(n22133)
         );
  NR2 U23943 ( .I1(n22172), .I2(n22118), .O(n22073) );
  NR2 U23944 ( .I1(n22166), .I2(n17195), .O(n22078) );
  NR2 U23945 ( .I1(n22169), .I2(n22121), .O(n22077) );
  INV1S U23946 ( .I(template_store[2]), .O(n22101) );
  NR2 U23947 ( .I1(n22101), .I2(n22168), .O(n22070) );
  NR2 U23948 ( .I1(n22170), .I2(n22162), .O(n22069) );
  HA1 U23949 ( .A(n22067), .B(n22066), .C(n22068), .S(n22063) );
  NR2 U23950 ( .I1(n22167), .I2(n13810), .O(n22081) );
  NR2 U23951 ( .I1(n22122), .I2(n22171), .O(n22080) );
  NR2 U23952 ( .I1(n22122), .I2(n22168), .O(n22141) );
  NR2 U23953 ( .I1(n22101), .I2(n13810), .O(n22140) );
  NR2 U23954 ( .I1(n22172), .I2(n17195), .O(n22100) );
  NR2 U23955 ( .I1(n22170), .I2(n22121), .O(n22099) );
  NR2 U23956 ( .I1(n22172), .I2(n22162), .O(n22098) );
  FA1S U23957 ( .A(n22070), .B(n22069), .CI(n22068), .CO(n22097), .S(n22075)
         );
  FA1S U23958 ( .A(n22073), .B(n22072), .CI(n22071), .CO(n22096), .S(n22076)
         );
  FA1S U23959 ( .A(n22076), .B(n22075), .CI(n22074), .CO(n22083), .S(n22151)
         );
  NR2 U23960 ( .I1(n22167), .I2(n22168), .O(n22095) );
  NR2 U23961 ( .I1(n22122), .I2(n13809), .O(n22094) );
  NR2 U23962 ( .I1(n22166), .I2(n22121), .O(n22089) );
  NR2 U23963 ( .I1(n22169), .I2(n22118), .O(n22088) );
  NR2 U23964 ( .I1(n22170), .I2(n13810), .O(n22087) );
  NR2 U23965 ( .I1(n22101), .I2(n22171), .O(n22086) );
  HA1 U23966 ( .A(n22078), .B(n22077), .C(n22085), .S(n22071) );
  FA1S U23967 ( .A(n22081), .B(n22080), .CI(n22079), .CO(n22090), .S(n22074)
         );
  NR2 U23968 ( .I1(n22156), .I2(n22157), .O(n22261) );
  FA1S U23969 ( .A(n22084), .B(n22083), .CI(n22082), .CO(n22158), .S(n22157)
         );
  NR2 U23970 ( .I1(n22172), .I2(n13810), .O(n22184) );
  FA1S U23971 ( .A(n22087), .B(n22086), .CI(n22085), .CO(n22183), .S(n22091)
         );
  NR2 U23972 ( .I1(n22166), .I2(n22118), .O(n22175) );
  NR2 U23973 ( .I1(n22101), .I2(n13809), .O(n22174) );
  FA1S U23974 ( .A(n22092), .B(n22091), .CI(n22090), .CO(n22192), .S(n22082)
         );
  NR2 U23975 ( .I1(n22170), .I2(n22168), .O(n22165) );
  NR2 U23976 ( .I1(n22169), .I2(n22162), .O(n22164) );
  NR2 U23977 ( .I1(n22167), .I2(n22171), .O(n22163) );
  FA1S U23978 ( .A(n22095), .B(n22094), .CI(n22093), .CO(n22189), .S(n22092)
         );
  FA1S U23979 ( .A(n22098), .B(n22097), .CI(n22096), .CO(n22188), .S(n22084)
         );
  NR2 U23980 ( .I1(n22158), .I2(n22159), .O(n22255) );
  NR2 U23981 ( .I1(n22261), .I2(n22255), .O(n22161) );
  NR2 U23982 ( .I1(n22293), .I2(n13810), .O(n22112) );
  NR2 U23983 ( .I1(n22167), .I2(n17195), .O(n22114) );
  NR2 U23984 ( .I1(n22101), .I2(n22121), .O(n22113) );
  NR2 U23985 ( .I1(n22122), .I2(n22118), .O(n22117) );
  NR2 U23986 ( .I1(n22293), .I2(n22162), .O(n22116) );
  NR2 U23987 ( .I1(n22101), .I2(n17195), .O(n22120) );
  NR2 U23988 ( .I1(n22122), .I2(n22121), .O(n22119) );
  NR2 U23989 ( .I1(n22167), .I2(n22118), .O(n22138) );
  NR2 U23990 ( .I1(n22101), .I2(n22162), .O(n22137) );
  HA1 U23991 ( .A(n22100), .B(n22099), .C(n22139), .S(n22136) );
  NR2 U23992 ( .I1(n22101), .I2(n22118), .O(n22109) );
  NR2 U23993 ( .I1(n22122), .I2(n22162), .O(n22108) );
  HA1 U23994 ( .A(n22103), .B(n22102), .C(n22104), .S(n22107) );
  FA1S U23995 ( .A(n22106), .B(n22105), .CI(n22104), .CO(n22134), .S(n22142)
         );
  NR2 U23996 ( .I1(n22131), .I2(n22132), .O(n22275) );
  FA1S U23997 ( .A(n22109), .B(n22108), .CI(n22107), .CO(n22143), .S(n22128)
         );
  FA1S U23998 ( .A(n22112), .B(n22111), .CI(n22110), .CO(n22131), .S(n22129)
         );
  OR2 U23999 ( .I1(n22128), .I2(n22129), .O(n22281) );
  FA1S U24000 ( .A(n22117), .B(n22116), .CI(n22115), .CO(n22110), .S(n22127)
         );
  NR2 U24001 ( .I1(n22126), .I2(n22127), .O(n22284) );
  NR2 U24002 ( .I1(n22293), .I2(n22118), .O(n22123) );
  NR2 U24003 ( .I1(n22293), .I2(n22121), .O(n22294) );
  NR2 U24004 ( .I1(n22122), .I2(n17195), .O(n22295) );
  ND2S U24005 ( .I1(n22294), .I2(n22295), .O(n22296) );
  INV1S U24006 ( .I(n22296), .O(n22292) );
  ND2S U24007 ( .I1(n22124), .I2(n22123), .O(n22289) );
  INV1S U24008 ( .I(n22289), .O(n22125) );
  AOI12HS U24009 ( .B1(n22290), .B2(n22292), .A1(n22125), .O(n22288) );
  OAI12HS U24010 ( .B1(n22284), .B2(n22288), .A1(n22285), .O(n22283) );
  INV1S U24011 ( .I(n22280), .O(n22130) );
  AOI12HS U24012 ( .B1(n22281), .B2(n22283), .A1(n22130), .O(n22279) );
  OAI12HS U24013 ( .B1(n22275), .B2(n22279), .A1(n22276), .O(n22274) );
  FA1S U24014 ( .A(n22135), .B(n22134), .CI(n22133), .CO(n22152), .S(n22145)
         );
  FA1S U24015 ( .A(n22138), .B(n22137), .CI(n22136), .CO(n22150), .S(n22144)
         );
  FA1S U24016 ( .A(n22141), .B(n22140), .CI(n22139), .CO(n22079), .S(n22149)
         );
  FA1S U24017 ( .A(n22144), .B(n22143), .CI(n22142), .CO(n22148), .S(n22132)
         );
  OR2 U24018 ( .I1(n22145), .I2(n22146), .O(n22272) );
  INV1S U24019 ( .I(n22271), .O(n22147) );
  AOI12HS U24020 ( .B1(n22274), .B2(n22272), .A1(n22147), .O(n22270) );
  FA1S U24021 ( .A(n22150), .B(n22149), .CI(n22148), .CO(n22154), .S(n22146)
         );
  FA1S U24022 ( .A(n22153), .B(n22152), .CI(n22151), .CO(n22156), .S(n22155)
         );
  NR2 U24023 ( .I1(n22154), .I2(n22155), .O(n22266) );
  OAI12HS U24024 ( .B1(n22270), .B2(n22266), .A1(n22267), .O(n22258) );
  ND2 U24025 ( .I1(n22157), .I2(n22156), .O(n22262) );
  ND2 U24026 ( .I1(n22159), .I2(n22158), .O(n22256) );
  OAI12HS U24027 ( .B1(n22255), .B2(n22262), .A1(n22256), .O(n22160) );
  AOI12H U24028 ( .B1(n22161), .B2(n22258), .A1(n22160), .O(n22246) );
  NR2 U24029 ( .I1(n22169), .I2(n13810), .O(n22181) );
  NR2 U24030 ( .I1(n22166), .I2(n22162), .O(n22180) );
  FA1S U24031 ( .A(n22165), .B(n22164), .CI(n22163), .CO(n22179), .S(n22190)
         );
  NR2 U24032 ( .I1(n22166), .I2(n13810), .O(n22208) );
  NR2 U24033 ( .I1(n22172), .I2(n22168), .O(n22178) );
  NR2 U24034 ( .I1(n22167), .I2(n13809), .O(n22177) );
  NR2 U24035 ( .I1(n22170), .I2(n22171), .O(n22176) );
  NR2 U24036 ( .I1(n22169), .I2(n22168), .O(n22202) );
  NR2 U24037 ( .I1(n22170), .I2(n13809), .O(n22201) );
  NR2 U24038 ( .I1(n22172), .I2(n22171), .O(n22200) );
  FA1S U24039 ( .A(n22175), .B(n22174), .CI(n22173), .CO(n22187), .S(n22182)
         );
  FA1S U24040 ( .A(n22178), .B(n22177), .CI(n22176), .CO(n22207), .S(n22186)
         );
  FA1S U24041 ( .A(n22181), .B(n22180), .CI(n22179), .CO(n22214), .S(n22185)
         );
  FA1S U24042 ( .A(n22184), .B(n22183), .CI(n22182), .CO(n22196), .S(n22193)
         );
  FA1S U24043 ( .A(n22187), .B(n22186), .CI(n22185), .CO(n22212), .S(n22195)
         );
  FA1S U24044 ( .A(n22190), .B(n22189), .CI(n22188), .CO(n22194), .S(n22191)
         );
  NR2 U24045 ( .I1(n22217), .I2(n22218), .O(n22243) );
  FA1S U24046 ( .A(n22193), .B(n22192), .CI(n22191), .CO(n22215), .S(n22159)
         );
  FA1S U24047 ( .A(n22196), .B(n22195), .CI(n22194), .CO(n22218), .S(n22216)
         );
  NR2 U24048 ( .I1(n22215), .I2(n22216), .O(n22247) );
  NR2 U24049 ( .I1(n22243), .I2(n22247), .O(n22231) );
  FA1S U24050 ( .A(n22199), .B(n22198), .CI(n22197), .CO(n22057), .S(n22221)
         );
  FA1S U24051 ( .A(n22202), .B(n22201), .CI(n22200), .CO(n22211), .S(n22206)
         );
  FA1S U24052 ( .A(n22205), .B(n22204), .CI(n22203), .CO(n22197), .S(n22210)
         );
  FA1S U24053 ( .A(n22208), .B(n22207), .CI(n22206), .CO(n22209), .S(n22213)
         );
  NR2 U24054 ( .I1(n22221), .I2(n22222), .O(n22228) );
  FA1S U24055 ( .A(n22211), .B(n22210), .CI(n22209), .CO(n22222), .S(n22219)
         );
  FA1S U24056 ( .A(n22214), .B(n22213), .CI(n22212), .CO(n22220), .S(n22217)
         );
  NR2 U24057 ( .I1(n22219), .I2(n22220), .O(n22235) );
  NR2 U24058 ( .I1(n22228), .I2(n22235), .O(n22224) );
  ND2 U24059 ( .I1(n22218), .I2(n22217), .O(n22244) );
  OAI12HS U24060 ( .B1(n22243), .B2(n22251), .A1(n22244), .O(n22232) );
  OAI12HS U24061 ( .B1(n22239), .B2(n22228), .A1(n22229), .O(n22223) );
  AOI12HS U24062 ( .B1(n22232), .B2(n22224), .A1(n22223), .O(n22225) );
  OAI12HS U24063 ( .B1(n22246), .B2(n22226), .A1(n22225), .O(n22301) );
  XNR2HS U24064 ( .I1(n22227), .I2(n22301), .O(PE_N142) );
  INV1S U24065 ( .I(n22228), .O(n22230) );
  ND2S U24066 ( .I1(n22230), .I2(n22229), .O(n22238) );
  INV1S U24067 ( .I(n22231), .O(n22234) );
  INV1S U24068 ( .I(n22232), .O(n22233) );
  OAI12HS U24069 ( .B1(n22246), .B2(n22234), .A1(n22233), .O(n22241) );
  INV1S U24070 ( .I(n22235), .O(n22240) );
  INV1S U24071 ( .I(n22239), .O(n22236) );
  AOI12HS U24072 ( .B1(n22241), .B2(n22240), .A1(n22236), .O(n22237) );
  XOR2HS U24073 ( .I1(n22238), .I2(n22237), .O(PE_N141) );
  ND2S U24074 ( .I1(n22240), .I2(n22239), .O(n22242) );
  XNR2HS U24075 ( .I1(n22242), .I2(n22241), .O(PE_N140) );
  INV1S U24076 ( .I(n22243), .O(n22245) );
  INV1S U24077 ( .I(n22247), .O(n22252) );
  INV1S U24078 ( .I(n22251), .O(n22248) );
  AOI12HS U24079 ( .B1(n22253), .B2(n22252), .A1(n22248), .O(n22249) );
  XOR2HS U24080 ( .I1(n22250), .I2(n22249), .O(PE_N139) );
  XNR2HS U24081 ( .I1(n22254), .I2(n22253), .O(PE_N138) );
  INV1S U24082 ( .I(n22255), .O(n22257) );
  INV1S U24083 ( .I(n22258), .O(n22265) );
  OAI12HS U24084 ( .B1(n22265), .B2(n22261), .A1(n22262), .O(n22259) );
  XNR2HS U24085 ( .I1(n22260), .I2(n22259), .O(PE_N137) );
  INV1S U24086 ( .I(n22261), .O(n22263) );
  XOR2HS U24087 ( .I1(n22265), .I2(n22264), .O(PE_N136) );
  INV1S U24088 ( .I(n22266), .O(n22268) );
  ND2S U24089 ( .I1(n22268), .I2(n22267), .O(n22269) );
  XOR2HS U24090 ( .I1(n22270), .I2(n22269), .O(PE_N135) );
  ND2S U24091 ( .I1(n22272), .I2(n22271), .O(n22273) );
  XNR2HS U24092 ( .I1(n22274), .I2(n22273), .O(PE_N134) );
  INV1S U24093 ( .I(n22275), .O(n22277) );
  ND2S U24094 ( .I1(n22277), .I2(n22276), .O(n22278) );
  XOR2HS U24095 ( .I1(n22279), .I2(n22278), .O(PE_N133) );
  ND2S U24096 ( .I1(n22281), .I2(n22280), .O(n22282) );
  XNR2HS U24097 ( .I1(n22283), .I2(n22282), .O(PE_N132) );
  INV1S U24098 ( .I(n22284), .O(n22286) );
  ND2S U24099 ( .I1(n22286), .I2(n22285), .O(n22287) );
  XOR2HS U24100 ( .I1(n22288), .I2(n22287), .O(PE_N131) );
  ND2S U24101 ( .I1(n22290), .I2(n22289), .O(n22291) );
  XNR2HS U24102 ( .I1(n22292), .I2(n22291), .O(PE_N130) );
  NR2 U24103 ( .I1(n22293), .I2(n17195), .O(PE_N128) );
  OR2S U24104 ( .I1(n22295), .I2(n22294), .O(n22297) );
  AN2S U24105 ( .I1(n22297), .I2(n22296), .O(PE_N129) );
  INV1S U24106 ( .I(n22298), .O(n22299) );
  AO12 U24107 ( .B1(n22301), .B2(n22300), .A1(n22299), .O(PE_N143) );
  NR2 U24108 ( .I1(n22332), .I2(n22324), .O(n22318) );
  NR2 U24109 ( .I1(n22332), .I2(n22302), .O(n22308) );
  NR2 U24110 ( .I1(n22348), .I2(n22324), .O(n22307) );
  FA1S U24111 ( .A(n22305), .B(n22304), .CI(n22303), .CO(n22306), .S(n22310)
         );
  FA1S U24112 ( .A(n22308), .B(n22307), .CI(n22306), .CO(n22317), .S(n22321)
         );
  FA1S U24113 ( .A(n22311), .B(n22310), .CI(n22309), .CO(n22320), .S(n22312)
         );
  NR2 U24114 ( .I1(n22312), .I2(n22313), .O(n22314) );
  MOAI1 U24115 ( .A1(n22315), .A2(n22314), .B1(n22313), .B2(n22312), .O(n22319) );
  FA1 U24116 ( .A(n22318), .B(n22317), .CI(n22316), .CO(PE_N95), .S(PE_N94) );
  FA1 U24117 ( .A(n22321), .B(n22320), .CI(n22319), .CO(n22316), .S(PE_N93) );
  NR2 U24118 ( .I1(n22332), .I2(n13813), .O(n22357) );
  NR2 U24119 ( .I1(n22323), .I2(n22322), .O(n22338) );
  NR2 U24120 ( .I1(n22325), .I2(n22324), .O(n22337) );
  HA1 U24121 ( .A(n22327), .B(n22326), .C(n22336), .S(n22352) );
  FA1S U24122 ( .A(n22330), .B(n22329), .CI(n22328), .CO(n21715), .S(n22355)
         );
  NR2 U24123 ( .I1(n22332), .I2(n22331), .O(n22347) );
  NR2 U24124 ( .I1(n22333), .I2(n13815), .O(n22346) );
  HA1 U24125 ( .A(n22335), .B(n22334), .C(n22342), .S(n22345) );
  FA1S U24126 ( .A(n22344), .B(n22343), .CI(n22342), .CO(n22359), .S(n22363)
         );
  NR2 U24127 ( .I1(n22348), .I2(n13813), .O(n22366) );
  FA1 U24128 ( .A(n22351), .B(n22350), .CI(n22349), .CO(n22365), .S(n22368) );
  FA1 U24129 ( .A(n22354), .B(n22353), .CI(n22352), .CO(n22364), .S(n22375) );
  FA1S U24130 ( .A(n22360), .B(n22359), .CI(n22358), .CO(n22405), .S(n22399)
         );
  NR2 U24131 ( .I1(n22401), .I2(n22402), .O(mult_x_433_n7) );
  FA1 U24132 ( .A(n22369), .B(n22368), .CI(n22367), .CO(n22395), .S(n22373) );
  ND2S U24133 ( .I1(n22404), .I2(n22403), .O(mult_x_433_n13) );
  NR2 U24134 ( .I1(n22403), .I2(n22404), .O(mult_x_433_n12) );
  FA1 U24135 ( .A(n22378), .B(n22377), .CI(n22376), .CO(mult_x_433_n14), .S(
        PE_N87) );
  FA1 U24136 ( .A(n22381), .B(n22380), .CI(n22379), .CO(n22376), .S(PE_N86) );
  FA1 U24137 ( .A(n22384), .B(n22383), .CI(n22382), .CO(n21722), .S(PE_N84) );
  FA1 U24138 ( .A(n22387), .B(n22386), .CI(n22385), .CO(n22382), .S(PE_N83) );
  FA1 U24139 ( .A(n22396), .B(n22395), .CI(n22394), .CO(mult_x_433_n51), .S(
        n22404) );
  NR2 U24140 ( .I1(n22397), .I2(n20735), .O(PE_N80) );
  FA1S U24141 ( .A(n22400), .B(n22399), .CI(n22398), .CO(mult_x_433_n33), .S(
        n22402) );
  FA1S U24142 ( .A(n22407), .B(n22406), .CI(n22405), .CO(n22313), .S(
        mult_x_433_n28) );
  HA1S U24143 ( .A(n22409), .B(n22408), .C(n22389), .S(PE_N81) );
  INV1S U24144 ( .I(template_store[23]), .O(n22527) );
  NR2 U24145 ( .I1(n22527), .I2(n22523), .O(n22413) );
  INV1S U24146 ( .I(template_store[22]), .O(n22529) );
  NR2 U24147 ( .I1(n22529), .I2(n22523), .O(n22557) );
  NR2 U24148 ( .I1(n22527), .I2(n13811), .O(n22556) );
  INV1S U24149 ( .I(template_store[21]), .O(n22530) );
  NR2 U24150 ( .I1(n22530), .I2(n22523), .O(n22563) );
  NR2 U24151 ( .I1(n22527), .I2(n22528), .O(n22562) );
  NR2 U24152 ( .I1(n22529), .I2(n13811), .O(n22561) );
  OR2S U24153 ( .I1(n22413), .I2(n22414), .O(n22659) );
  ND2S U24154 ( .I1(n22414), .I2(n22413), .O(n22657) );
  ND2S U24155 ( .I1(n22659), .I2(n22657), .O(n22585) );
  INV2 U24156 ( .I(n22415), .O(n22524) );
  NR2 U24157 ( .I1(n22530), .I2(n22524), .O(n22435) );
  INV1S U24158 ( .I(template_store[19]), .O(n22519) );
  NR2 U24159 ( .I1(n22519), .I2(n22528), .O(n22434) );
  NR2 U24160 ( .I1(n22530), .I2(n22461), .O(n22424) );
  INV1S U24161 ( .I(template_store[17]), .O(n22478) );
  NR2 U24162 ( .I1(n22478), .I2(n13811), .O(n22423) );
  NR2 U24163 ( .I1(n22529), .I2(n22479), .O(n22422) );
  NR2 U24164 ( .I1(n22529), .I2(n22461), .O(n22438) );
  NR2 U24165 ( .I1(n22478), .I2(n22523), .O(n22437) );
  INV1S U24166 ( .I(template_store[18]), .O(n22475) );
  NR2 U24167 ( .I1(n22475), .I2(n13811), .O(n22436) );
  INV2 U24168 ( .I(n22418), .O(n22526) );
  NR2 U24169 ( .I1(n22519), .I2(n22526), .O(n22444) );
  NR2 U24170 ( .I1(n22527), .I2(n22651), .O(n22443) );
  NR2 U24171 ( .I1(n22475), .I2(n22526), .O(n22446) );
  NR2 U24172 ( .I1(n22478), .I2(n22528), .O(n22445) );
  INV1S U24173 ( .I(template_store[20]), .O(n22525) );
  NR2 U24174 ( .I1(n22525), .I2(n22526), .O(n22441) );
  NR2 U24175 ( .I1(n22527), .I2(n22479), .O(n22440) );
  NR2 U24176 ( .I1(n22525), .I2(n22524), .O(n22421) );
  INV1S U24177 ( .I(template_store[16]), .O(n22652) );
  NR2 U24178 ( .I1(n22652), .I2(n22523), .O(n22427) );
  HA1 U24179 ( .A(n22421), .B(n22420), .C(n22439), .S(n22426) );
  NR2 U24180 ( .I1(n22525), .I2(n22461), .O(n22449) );
  NR2 U24181 ( .I1(n22652), .I2(n13811), .O(n22448) );
  NR2 U24182 ( .I1(n22530), .I2(n22479), .O(n22447) );
  NR2 U24183 ( .I1(n22519), .I2(n22524), .O(n22495) );
  NR2 U24184 ( .I1(n22529), .I2(n22651), .O(n22494) );
  NR2 U24185 ( .I1(n22478), .I2(n22526), .O(n22463) );
  NR2 U24186 ( .I1(n22652), .I2(n22528), .O(n22462) );
  FA1S U24187 ( .A(n22424), .B(n22423), .CI(n22422), .CO(n22429), .S(n22451)
         );
  FA1S U24188 ( .A(n22427), .B(n22426), .CI(n22425), .CO(n22431), .S(n22450)
         );
  FA1S U24189 ( .A(n22430), .B(n22429), .CI(n22428), .CO(n22551), .S(n22455)
         );
  FA1S U24190 ( .A(n22433), .B(n22432), .CI(n22431), .CO(n22550), .S(n22454)
         );
  NR2 U24191 ( .I1(n22530), .I2(n22526), .O(n22522) );
  NR2 U24192 ( .I1(n22475), .I2(n22523), .O(n22521) );
  NR2 U24193 ( .I1(n22519), .I2(n13811), .O(n22520) );
  NR2 U24194 ( .I1(n22529), .I2(n22524), .O(n22533) );
  NR2 U24195 ( .I1(n22525), .I2(n22528), .O(n22532) );
  NR2 U24196 ( .I1(n22527), .I2(n22461), .O(n22542) );
  FA1S U24197 ( .A(n22438), .B(n22437), .CI(n22436), .CO(n22541), .S(n22428)
         );
  FA1S U24198 ( .A(n22441), .B(n22440), .CI(n22439), .CO(n22540), .S(n22432)
         );
  NR2 U24199 ( .I1(n22515), .I2(n22516), .O(n22613) );
  FA1S U24200 ( .A(n22444), .B(n22443), .CI(n22442), .CO(n22433), .S(n22510)
         );
  NR2 U24201 ( .I1(n22475), .I2(n22524), .O(n22460) );
  NR2 U24202 ( .I1(n22530), .I2(n22651), .O(n22459) );
  NR2 U24203 ( .I1(n22652), .I2(n22526), .O(n22457) );
  NR2 U24204 ( .I1(n22475), .I2(n22461), .O(n22456) );
  FA1S U24205 ( .A(n22449), .B(n22448), .CI(n22447), .CO(n22425), .S(n22490)
         );
  FA1S U24206 ( .A(n22452), .B(n22451), .CI(n22450), .CO(n22453), .S(n22508)
         );
  FA1S U24207 ( .A(n22455), .B(n22454), .CI(n22453), .CO(n22515), .S(n22514)
         );
  NR2 U24208 ( .I1(n22513), .I2(n22514), .O(n22619) );
  NR2 U24209 ( .I1(n22613), .I2(n22619), .O(n22518) );
  NR2 U24210 ( .I1(n22519), .I2(n22479), .O(n22469) );
  NR2 U24211 ( .I1(n22475), .I2(n22479), .O(n22474) );
  NR2 U24212 ( .I1(n22519), .I2(n22651), .O(n22473) );
  NR2 U24213 ( .I1(n22652), .I2(n22461), .O(n22477) );
  NR2 U24214 ( .I1(n22478), .I2(n22479), .O(n22476) );
  NR2 U24215 ( .I1(n22478), .I2(n22524), .O(n22466) );
  NR2 U24216 ( .I1(n22525), .I2(n22651), .O(n22465) );
  NR2 U24217 ( .I1(n22652), .I2(n22524), .O(n22471) );
  NR2 U24218 ( .I1(n22478), .I2(n22461), .O(n22470) );
  FA1S U24219 ( .A(n22460), .B(n22459), .CI(n22458), .CO(n22491), .S(n22500)
         );
  NR2 U24220 ( .I1(n22519), .I2(n22461), .O(n22498) );
  NR2 U24221 ( .I1(n22525), .I2(n22479), .O(n22497) );
  NR2 U24222 ( .I1(n22488), .I2(n22489), .O(n22633) );
  FA1S U24223 ( .A(n22466), .B(n22465), .CI(n22464), .CO(n22501), .S(n22485)
         );
  FA1S U24224 ( .A(n22469), .B(n22468), .CI(n22467), .CO(n22488), .S(n22486)
         );
  OR2 U24225 ( .I1(n22485), .I2(n22486), .O(n22639) );
  FA1S U24226 ( .A(n22474), .B(n22473), .CI(n22472), .CO(n22467), .S(n22484)
         );
  NR2 U24227 ( .I1(n22483), .I2(n22484), .O(n22642) );
  NR2 U24228 ( .I1(n22475), .I2(n22651), .O(n22480) );
  NR2 U24229 ( .I1(n22478), .I2(n22651), .O(n22653) );
  NR2 U24230 ( .I1(n22652), .I2(n22479), .O(n22654) );
  ND2S U24231 ( .I1(n22653), .I2(n22654), .O(n22655) );
  INV1S U24232 ( .I(n22655), .O(n22650) );
  ND2S U24233 ( .I1(n22481), .I2(n22480), .O(n22647) );
  INV1S U24234 ( .I(n22647), .O(n22482) );
  AOI12HS U24235 ( .B1(n22648), .B2(n22650), .A1(n22482), .O(n22646) );
  OAI12HS U24236 ( .B1(n22642), .B2(n22646), .A1(n22643), .O(n22641) );
  INV1S U24237 ( .I(n22638), .O(n22487) );
  AOI12HS U24238 ( .B1(n22639), .B2(n22641), .A1(n22487), .O(n22637) );
  OAI12HS U24239 ( .B1(n22633), .B2(n22637), .A1(n22634), .O(n22632) );
  FA1S U24240 ( .A(n22492), .B(n22491), .CI(n22490), .CO(n22509), .S(n22502)
         );
  FA1S U24241 ( .A(n22495), .B(n22494), .CI(n22493), .CO(n22452), .S(n22507)
         );
  FA1S U24242 ( .A(n22498), .B(n22497), .CI(n22496), .CO(n22506), .S(n22499)
         );
  FA1S U24243 ( .A(n22501), .B(n22500), .CI(n22499), .CO(n22505), .S(n22489)
         );
  OR2 U24244 ( .I1(n22502), .I2(n22503), .O(n22630) );
  INV1S U24245 ( .I(n22629), .O(n22504) );
  AOI12HS U24246 ( .B1(n22632), .B2(n22630), .A1(n22504), .O(n22628) );
  FA1S U24247 ( .A(n22507), .B(n22506), .CI(n22505), .CO(n22511), .S(n22503)
         );
  FA1S U24248 ( .A(n22510), .B(n22509), .CI(n22508), .CO(n22513), .S(n22512)
         );
  NR2 U24249 ( .I1(n22511), .I2(n22512), .O(n22624) );
  ND2 U24250 ( .I1(n22514), .I2(n22513), .O(n22620) );
  OAI12HS U24251 ( .B1(n22620), .B2(n22613), .A1(n22614), .O(n22517) );
  AOI12H U24252 ( .B1(n22518), .B2(n22616), .A1(n22517), .O(n22604) );
  NR2 U24253 ( .I1(n22529), .I2(n22526), .O(n22539) );
  NR2 U24254 ( .I1(n22519), .I2(n22523), .O(n22538) );
  FA1S U24255 ( .A(n22522), .B(n22521), .CI(n22520), .CO(n22537), .S(n22548)
         );
  NR2 U24256 ( .I1(n22525), .I2(n22523), .O(n22566) );
  NR2 U24257 ( .I1(n22527), .I2(n22524), .O(n22536) );
  NR2 U24258 ( .I1(n22530), .I2(n22528), .O(n22535) );
  NR2 U24259 ( .I1(n22525), .I2(n13811), .O(n22534) );
  NR2 U24260 ( .I1(n22527), .I2(n22526), .O(n22560) );
  NR2 U24261 ( .I1(n22529), .I2(n22528), .O(n22559) );
  NR2 U24262 ( .I1(n22530), .I2(n13811), .O(n22558) );
  FA1S U24263 ( .A(n22533), .B(n22532), .CI(n22531), .CO(n22545), .S(n22547)
         );
  FA1S U24264 ( .A(n22536), .B(n22535), .CI(n22534), .CO(n22565), .S(n22544)
         );
  FA1S U24265 ( .A(n22539), .B(n22538), .CI(n22537), .CO(n22572), .S(n22543)
         );
  FA1S U24266 ( .A(n22542), .B(n22541), .CI(n22540), .CO(n22554), .S(n22546)
         );
  FA1S U24267 ( .A(n22545), .B(n22544), .CI(n22543), .CO(n22570), .S(n22553)
         );
  FA1S U24268 ( .A(n22548), .B(n22547), .CI(n22546), .CO(n22552), .S(n22549)
         );
  NR2 U24269 ( .I1(n22575), .I2(n22576), .O(n22601) );
  FA1S U24270 ( .A(n22551), .B(n22550), .CI(n22549), .CO(n22573), .S(n22516)
         );
  FA1S U24271 ( .A(n22554), .B(n22553), .CI(n22552), .CO(n22576), .S(n22574)
         );
  NR2 U24272 ( .I1(n22573), .I2(n22574), .O(n22605) );
  NR2 U24273 ( .I1(n22601), .I2(n22605), .O(n22589) );
  FA1S U24274 ( .A(n22557), .B(n22556), .CI(n22555), .CO(n22414), .S(n22579)
         );
  FA1S U24275 ( .A(n22560), .B(n22559), .CI(n22558), .CO(n22569), .S(n22564)
         );
  FA1S U24276 ( .A(n22563), .B(n22562), .CI(n22561), .CO(n22555), .S(n22568)
         );
  FA1S U24277 ( .A(n22566), .B(n22565), .CI(n22564), .CO(n22567), .S(n22571)
         );
  NR2 U24278 ( .I1(n22579), .I2(n22580), .O(n22586) );
  FA1S U24279 ( .A(n22569), .B(n22568), .CI(n22567), .CO(n22580), .S(n22577)
         );
  FA1S U24280 ( .A(n22572), .B(n22571), .CI(n22570), .CO(n22578), .S(n22575)
         );
  NR2 U24281 ( .I1(n22577), .I2(n22578), .O(n22593) );
  NR2 U24282 ( .I1(n22586), .I2(n22593), .O(n22582) );
  ND2 U24283 ( .I1(n22574), .I2(n22573), .O(n22609) );
  ND2 U24284 ( .I1(n22576), .I2(n22575), .O(n22602) );
  OAI12HS U24285 ( .B1(n22609), .B2(n22601), .A1(n22602), .O(n22590) );
  OAI12HS U24286 ( .B1(n22597), .B2(n22586), .A1(n22587), .O(n22581) );
  AOI12HS U24287 ( .B1(n22590), .B2(n22582), .A1(n22581), .O(n22583) );
  OAI12HS U24288 ( .B1(n22604), .B2(n22584), .A1(n22583), .O(n22660) );
  XNR2HS U24289 ( .I1(n22585), .I2(n22660), .O(PE_N110) );
  INV1S U24290 ( .I(n22586), .O(n22588) );
  ND2S U24291 ( .I1(n22588), .I2(n22587), .O(n22596) );
  INV1S U24292 ( .I(n22589), .O(n22592) );
  INV1S U24293 ( .I(n22590), .O(n22591) );
  INV1S U24294 ( .I(n22593), .O(n22598) );
  INV1S U24295 ( .I(n22597), .O(n22594) );
  XOR2HS U24296 ( .I1(n22596), .I2(n22595), .O(PE_N109) );
  ND2S U24297 ( .I1(n22598), .I2(n22597), .O(n22600) );
  XNR2HS U24298 ( .I1(n22600), .I2(n22599), .O(PE_N108) );
  INV1S U24299 ( .I(n22601), .O(n22603) );
  INV1 U24300 ( .I(n22604), .O(n22611) );
  INV1S U24301 ( .I(n22605), .O(n22610) );
  INV1S U24302 ( .I(n22609), .O(n22606) );
  AOI12HS U24303 ( .B1(n22611), .B2(n22610), .A1(n22606), .O(n22607) );
  XOR2HS U24304 ( .I1(n22608), .I2(n22607), .O(PE_N107) );
  XNR2HS U24305 ( .I1(n22612), .I2(n22611), .O(PE_N106) );
  INV1S U24306 ( .I(n22613), .O(n22615) );
  INV1S U24307 ( .I(n22616), .O(n22623) );
  OAI12HS U24308 ( .B1(n22623), .B2(n22619), .A1(n22620), .O(n22617) );
  XNR2HS U24309 ( .I1(n22618), .I2(n22617), .O(PE_N105) );
  INV1S U24310 ( .I(n22619), .O(n22621) );
  XOR2HS U24311 ( .I1(n22623), .I2(n22622), .O(PE_N104) );
  INV1S U24312 ( .I(n22624), .O(n22626) );
  XOR2HS U24313 ( .I1(n22628), .I2(n22627), .O(PE_N103) );
  ND2S U24314 ( .I1(n22630), .I2(n22629), .O(n22631) );
  XNR2HS U24315 ( .I1(n22632), .I2(n22631), .O(PE_N102) );
  INV1S U24316 ( .I(n22633), .O(n22635) );
  ND2S U24317 ( .I1(n22635), .I2(n22634), .O(n22636) );
  XOR2HS U24318 ( .I1(n22637), .I2(n22636), .O(PE_N101) );
  ND2S U24319 ( .I1(n22639), .I2(n22638), .O(n22640) );
  XNR2HS U24320 ( .I1(n22641), .I2(n22640), .O(PE_N100) );
  INV1S U24321 ( .I(n22642), .O(n22644) );
  ND2S U24322 ( .I1(n22644), .I2(n22643), .O(n22645) );
  XOR2HS U24323 ( .I1(n22646), .I2(n22645), .O(PE_N99) );
  ND2S U24324 ( .I1(n22648), .I2(n22647), .O(n22649) );
  XNR2HS U24325 ( .I1(n22650), .I2(n22649), .O(PE_N98) );
  NR2 U24326 ( .I1(n22652), .I2(n22651), .O(PE_N96) );
  OR2S U24327 ( .I1(n22654), .I2(n22653), .O(n22656) );
  AN2S U24328 ( .I1(n22656), .I2(n22655), .O(PE_N97) );
  INV1S U24329 ( .I(n22657), .O(n22658) );
  AO12 U24330 ( .B1(n22660), .B2(n22659), .A1(n22658), .O(PE_N111) );
  INV1S U24331 ( .I(template_store[63]), .O(n22777) );
  NR2 U24332 ( .I1(n22777), .I2(n22778), .O(n22664) );
  NR2 U24333 ( .I1(n22777), .I2(n22773), .O(n22825) );
  INV1S U24334 ( .I(template_store[62]), .O(n22780) );
  NR2 U24335 ( .I1(n22780), .I2(n22778), .O(n22824) );
  NR2 U24336 ( .I1(n22780), .I2(n22773), .O(n22816) );
  INV1S U24337 ( .I(template_store[61]), .O(n22775) );
  NR2 U24338 ( .I1(n22775), .I2(n22778), .O(n22815) );
  NR2 U24339 ( .I1(n22777), .I2(n20728), .O(n22814) );
  NR2 U24340 ( .I1(n22664), .I2(n22665), .O(n22841) );
  INV1S U24341 ( .I(n22841), .O(n22666) );
  ND2S U24342 ( .I1(n22665), .I2(n22664), .O(n22840) );
  ND2S U24343 ( .I1(n22666), .I2(n22840), .O(n22837) );
  NR2 U24344 ( .I1(n22775), .I2(n22713), .O(n22679) );
  NR2 U24345 ( .I1(n22780), .I2(n22730), .O(n22678) );
  INV1S U24346 ( .I(template_store[58]), .O(n22714) );
  NR2 U24347 ( .I1(n22714), .I2(n22776), .O(n22673) );
  INV1S U24348 ( .I(template_store[56]), .O(n22910) );
  NR2 U24349 ( .I1(n22910), .I2(n22773), .O(n22672) );
  NR2 U24350 ( .I1(n22780), .I2(n22909), .O(n22742) );
  NR2 U24351 ( .I1(n22775), .I2(n22909), .O(n22712) );
  INV1S U24352 ( .I(template_store[60]), .O(n22779) );
  NR2 U24353 ( .I1(n22779), .I2(n22730), .O(n22711) );
  NR2 U24354 ( .I1(n22910), .I2(n22776), .O(n22716) );
  INV1S U24355 ( .I(template_store[57]), .O(n22731) );
  INV2 U24356 ( .I(n22671), .O(n22769) );
  NR2 U24357 ( .I1(n22731), .I2(n22769), .O(n22715) );
  INV1S U24358 ( .I(template_store[59]), .O(n22774) );
  NR2 U24359 ( .I1(n22774), .I2(n22769), .O(n22676) );
  NR2 U24360 ( .I1(n22775), .I2(n22730), .O(n22675) );
  NR2 U24361 ( .I1(n22731), .I2(n22776), .O(n22709) );
  NR2 U24362 ( .I1(n22714), .I2(n22769), .O(n22708) );
  NR2 U24363 ( .I1(n22779), .I2(n22713), .O(n22745) );
  NR2 U24364 ( .I1(n22731), .I2(n20728), .O(n22744) );
  NR2 U24365 ( .I1(n22779), .I2(n22769), .O(n22682) );
  NR2 U24366 ( .I1(n22714), .I2(n20728), .O(n22681) );
  NR2 U24367 ( .I1(n22774), .I2(n22776), .O(n22687) );
  NR2 U24368 ( .I1(n22731), .I2(n22773), .O(n22686) );
  NR2 U24369 ( .I1(n22910), .I2(n22778), .O(n22690) );
  NR2 U24370 ( .I1(n22777), .I2(n22909), .O(n22689) );
  FA1S U24371 ( .A(n22676), .B(n22675), .CI(n22674), .CO(n22688), .S(n22740)
         );
  NR2 U24372 ( .I1(n22731), .I2(n22778), .O(n22707) );
  FA1S U24373 ( .A(n22679), .B(n22678), .CI(n22677), .CO(n22706), .S(n22760)
         );
  FA1S U24374 ( .A(n22682), .B(n22681), .CI(n22680), .CO(n22705), .S(n22684)
         );
  FA1S U24375 ( .A(n22685), .B(n22684), .CI(n22683), .CO(n22692), .S(n22758)
         );
  NR2 U24376 ( .I1(n22775), .I2(n22769), .O(n22696) );
  NR2 U24377 ( .I1(n22777), .I2(n22730), .O(n22695) );
  NR2 U24378 ( .I1(n22780), .I2(n22713), .O(n22704) );
  NR2 U24379 ( .I1(n22774), .I2(n20728), .O(n22703) );
  NR2 U24380 ( .I1(n22779), .I2(n22776), .O(n22698) );
  NR2 U24381 ( .I1(n22714), .I2(n22773), .O(n22697) );
  FA1S U24382 ( .A(n22690), .B(n22689), .CI(n22688), .CO(n22699), .S(n22683)
         );
  NR2 U24383 ( .I1(n22763), .I2(n22764), .O(n22875) );
  FA1S U24384 ( .A(n22693), .B(n22692), .CI(n22691), .CO(n22765), .S(n22764)
         );
  NR2 U24385 ( .I1(n22780), .I2(n22769), .O(n22792) );
  FA1S U24386 ( .A(n22696), .B(n22695), .CI(n22694), .CO(n22791), .S(n22701)
         );
  NR2 U24387 ( .I1(n22775), .I2(n22776), .O(n22783) );
  NR2 U24388 ( .I1(n22779), .I2(n20728), .O(n22782) );
  FA1S U24389 ( .A(n22701), .B(n22700), .CI(n22699), .CO(n22800), .S(n22691)
         );
  NR2 U24390 ( .I1(n22774), .I2(n22773), .O(n22772) );
  NR2 U24391 ( .I1(n22777), .I2(n22713), .O(n22771) );
  NR2 U24392 ( .I1(n22714), .I2(n22778), .O(n22770) );
  FA1S U24393 ( .A(n22704), .B(n22703), .CI(n22702), .CO(n22797), .S(n22700)
         );
  FA1S U24394 ( .A(n22707), .B(n22706), .CI(n22705), .CO(n22796), .S(n22693)
         );
  NR2 U24395 ( .I1(n22765), .I2(n22766), .O(n22869) );
  NR2 U24396 ( .I1(n22875), .I2(n22869), .O(n22768) );
  NR2 U24397 ( .I1(n22779), .I2(n22909), .O(n22722) );
  NR2 U24398 ( .I1(n22731), .I2(n22713), .O(n22724) );
  NR2 U24399 ( .I1(n22714), .I2(n22730), .O(n22723) );
  NR2 U24400 ( .I1(n22910), .I2(n22769), .O(n22727) );
  NR2 U24401 ( .I1(n22774), .I2(n22909), .O(n22726) );
  NR2 U24402 ( .I1(n22910), .I2(n22713), .O(n22729) );
  NR2 U24403 ( .I1(n22714), .I2(n22909), .O(n22728) );
  NR2 U24404 ( .I1(n22774), .I2(n22713), .O(n22748) );
  NR2 U24405 ( .I1(n22910), .I2(n20728), .O(n22747) );
  FA1S U24406 ( .A(n22712), .B(n22711), .CI(n22710), .CO(n22741), .S(n22750)
         );
  NR2 U24407 ( .I1(n22714), .I2(n22713), .O(n22719) );
  NR2 U24408 ( .I1(n22774), .I2(n22730), .O(n22718) );
  NR2 U24409 ( .I1(n22738), .I2(n22739), .O(n22889) );
  FA1S U24410 ( .A(n22719), .B(n22718), .CI(n22717), .CO(n22749), .S(n22735)
         );
  FA1S U24411 ( .A(n22722), .B(n22721), .CI(n22720), .CO(n22738), .S(n22736)
         );
  FA1S U24412 ( .A(n22727), .B(n22726), .CI(n22725), .CO(n22720), .S(n22734)
         );
  NR2 U24413 ( .I1(n22733), .I2(n22734), .O(n22898) );
  NR2 U24414 ( .I1(n22910), .I2(n22730), .O(n22911) );
  NR2 U24415 ( .I1(n22731), .I2(n22909), .O(n22912) );
  ND2S U24416 ( .I1(n22911), .I2(n22912), .O(n22913) );
  INV1S U24417 ( .I(n22913), .O(n22908) );
  NR2 U24418 ( .I1(n22731), .I2(n22730), .O(n22904) );
  ND2S U24419 ( .I1(n22903), .I2(n22904), .O(n22905) );
  INV1S U24420 ( .I(n22905), .O(n22732) );
  NR2 U24421 ( .I1(n22908), .I2(n22732), .O(n22902) );
  ND2S U24422 ( .I1(n22734), .I2(n22733), .O(n22899) );
  OAI12HS U24423 ( .B1(n22898), .B2(n22902), .A1(n22899), .O(n22897) );
  INV1S U24424 ( .I(n22894), .O(n22737) );
  AOI12HS U24425 ( .B1(n22895), .B2(n22897), .A1(n22737), .O(n22893) );
  OAI12HS U24426 ( .B1(n22889), .B2(n22893), .A1(n22890), .O(n22887) );
  FA1S U24427 ( .A(n22742), .B(n22741), .CI(n22740), .CO(n22759), .S(n22752)
         );
  FA1S U24428 ( .A(n22745), .B(n22744), .CI(n22743), .CO(n22685), .S(n22757)
         );
  FA1S U24429 ( .A(n22748), .B(n22747), .CI(n22746), .CO(n22756), .S(n22751)
         );
  FA1S U24430 ( .A(n22751), .B(n22750), .CI(n22749), .CO(n22755), .S(n22739)
         );
  OR2 U24431 ( .I1(n22752), .I2(n22753), .O(n22886) );
  INV1S U24432 ( .I(n22885), .O(n22754) );
  AOI12HS U24433 ( .B1(n22887), .B2(n22886), .A1(n22754), .O(n22884) );
  FA1S U24434 ( .A(n22757), .B(n22756), .CI(n22755), .CO(n22761), .S(n22753)
         );
  FA1S U24435 ( .A(n22760), .B(n22759), .CI(n22758), .CO(n22763), .S(n22762)
         );
  NR2 U24436 ( .I1(n22761), .I2(n22762), .O(n22880) );
  OAI12HS U24437 ( .B1(n22884), .B2(n22880), .A1(n22881), .O(n22872) );
  ND2 U24438 ( .I1(n22764), .I2(n22763), .O(n22876) );
  OAI12HS U24439 ( .B1(n22869), .B2(n22876), .A1(n22870), .O(n22767) );
  NR2 U24440 ( .I1(n22779), .I2(n22773), .O(n22789) );
  NR2 U24441 ( .I1(n22777), .I2(n22769), .O(n22788) );
  FA1S U24442 ( .A(n22772), .B(n22771), .CI(n22770), .CO(n22787), .S(n22798)
         );
  NR2 U24443 ( .I1(n22775), .I2(n22773), .O(n22819) );
  NR2 U24444 ( .I1(n22780), .I2(n22776), .O(n22786) );
  NR2 U24445 ( .I1(n22774), .I2(n22778), .O(n22785) );
  NR2 U24446 ( .I1(n22775), .I2(n20728), .O(n22784) );
  NR2 U24447 ( .I1(n22777), .I2(n22776), .O(n22813) );
  NR2 U24448 ( .I1(n22779), .I2(n22778), .O(n22812) );
  NR2 U24449 ( .I1(n22780), .I2(n20728), .O(n22811) );
  FA1S U24450 ( .A(n22783), .B(n22782), .CI(n22781), .CO(n22795), .S(n22790)
         );
  FA1S U24451 ( .A(n22786), .B(n22785), .CI(n22784), .CO(n22818), .S(n22794)
         );
  FA1S U24452 ( .A(n22789), .B(n22788), .CI(n22787), .CO(n22822), .S(n22793)
         );
  FA1S U24453 ( .A(n22792), .B(n22791), .CI(n22790), .CO(n22804), .S(n22801)
         );
  FA1S U24454 ( .A(n22795), .B(n22794), .CI(n22793), .CO(n22820), .S(n22803)
         );
  FA1S U24455 ( .A(n22798), .B(n22797), .CI(n22796), .CO(n22802), .S(n22799)
         );
  NR2 U24456 ( .I1(n22807), .I2(n22808), .O(n22857) );
  FA1S U24457 ( .A(n22801), .B(n22800), .CI(n22799), .CO(n22805), .S(n22766)
         );
  FA1S U24458 ( .A(n22804), .B(n22803), .CI(n22802), .CO(n22808), .S(n22806)
         );
  NR2 U24459 ( .I1(n22805), .I2(n22806), .O(n22861) );
  NR2 U24460 ( .I1(n22857), .I2(n22861), .O(n22839) );
  INV1S U24461 ( .I(n22839), .O(n22810) );
  OAI12HS U24462 ( .B1(n22857), .B2(n22865), .A1(n22858), .O(n22845) );
  INV1S U24463 ( .I(n22845), .O(n22809) );
  FA1S U24464 ( .A(n22813), .B(n22812), .CI(n22811), .CO(n22828), .S(n22817)
         );
  FA1S U24465 ( .A(n22816), .B(n22815), .CI(n22814), .CO(n22823), .S(n22827)
         );
  FA1S U24466 ( .A(n22819), .B(n22818), .CI(n22817), .CO(n22826), .S(n22821)
         );
  FA1S U24467 ( .A(n22822), .B(n22821), .CI(n22820), .CO(n22830), .S(n22807)
         );
  FA1S U24468 ( .A(n22825), .B(n22824), .CI(n22823), .CO(n22665), .S(n22831)
         );
  FA1S U24469 ( .A(n22828), .B(n22827), .CI(n22826), .CO(n22832), .S(n22829)
         );
  ND2S U24470 ( .I1(n22854), .I2(n22849), .O(n22838) );
  INV1S U24471 ( .I(n22838), .O(n22835) );
  INV1S U24472 ( .I(n22853), .O(n22850) );
  ND2S U24473 ( .I1(n22832), .I2(n22831), .O(n22848) );
  INV1S U24474 ( .I(n22848), .O(n22833) );
  AOI12HS U24475 ( .B1(n22850), .B2(n22849), .A1(n22833), .O(n22842) );
  INV1S U24476 ( .I(n22842), .O(n22834) );
  AOI12HS U24477 ( .B1(n22855), .B2(n22835), .A1(n22834), .O(n22836) );
  XOR2HS U24478 ( .I1(n22837), .I2(n22836), .O(PE_N30) );
  NR2 U24479 ( .I1(n22841), .I2(n22838), .O(n22844) );
  ND2S U24480 ( .I1(n22839), .I2(n22844), .O(n22847) );
  OAI12HS U24481 ( .B1(n22842), .B2(n22841), .A1(n22840), .O(n22843) );
  AOI12HS U24482 ( .B1(n22845), .B2(n22844), .A1(n22843), .O(n22846) );
  OAI12HS U24483 ( .B1(n22860), .B2(n22847), .A1(n22846), .O(PE_N31) );
  ND2S U24484 ( .I1(n22849), .I2(n22848), .O(n22852) );
  AOI12HS U24485 ( .B1(n22855), .B2(n22854), .A1(n22850), .O(n22851) );
  XOR2HS U24486 ( .I1(n22852), .I2(n22851), .O(PE_N29) );
  ND2S U24487 ( .I1(n22854), .I2(n22853), .O(n22856) );
  XNR2HS U24488 ( .I1(n22856), .I2(n22855), .O(PE_N28) );
  INV1S U24489 ( .I(n22857), .O(n22859) );
  ND2S U24490 ( .I1(n22859), .I2(n22858), .O(n22864) );
  INV1S U24491 ( .I(n22861), .O(n22866) );
  INV1S U24492 ( .I(n22865), .O(n22862) );
  AOI12HS U24493 ( .B1(n22867), .B2(n22866), .A1(n22862), .O(n22863) );
  XOR2HS U24494 ( .I1(n22864), .I2(n22863), .O(PE_N27) );
  ND2S U24495 ( .I1(n22866), .I2(n22865), .O(n22868) );
  XNR2HS U24496 ( .I1(n22868), .I2(n22867), .O(PE_N26) );
  INV1S U24497 ( .I(n22869), .O(n22871) );
  ND2S U24498 ( .I1(n22871), .I2(n22870), .O(n22874) );
  INV1S U24499 ( .I(n22872), .O(n22879) );
  OAI12HS U24500 ( .B1(n22879), .B2(n22875), .A1(n22876), .O(n22873) );
  XNR2HS U24501 ( .I1(n22874), .I2(n22873), .O(PE_N25) );
  INV1S U24502 ( .I(n22875), .O(n22877) );
  ND2S U24503 ( .I1(n22877), .I2(n22876), .O(n22878) );
  XOR2HS U24504 ( .I1(n22879), .I2(n22878), .O(PE_N24) );
  INV1S U24505 ( .I(n22880), .O(n22882) );
  ND2S U24506 ( .I1(n22882), .I2(n22881), .O(n22883) );
  XOR2HS U24507 ( .I1(n22884), .I2(n22883), .O(PE_N23) );
  ND2S U24508 ( .I1(n22886), .I2(n22885), .O(n22888) );
  XNR2HS U24509 ( .I1(n22888), .I2(n22887), .O(PE_N22) );
  INV1S U24510 ( .I(n22889), .O(n22891) );
  ND2S U24511 ( .I1(n22891), .I2(n22890), .O(n22892) );
  XOR2HS U24512 ( .I1(n22893), .I2(n22892), .O(PE_N21) );
  ND2S U24513 ( .I1(n22895), .I2(n22894), .O(n22896) );
  XNR2HS U24514 ( .I1(n22897), .I2(n22896), .O(PE_N20) );
  INV1S U24515 ( .I(n22898), .O(n22900) );
  ND2S U24516 ( .I1(n22900), .I2(n22899), .O(n22901) );
  XOR2HS U24517 ( .I1(n22902), .I2(n22901), .O(PE_N19) );
  OR2S U24518 ( .I1(n22904), .I2(n22903), .O(n22906) );
  ND2S U24519 ( .I1(n22906), .I2(n22905), .O(n22907) );
  XNR2HS U24520 ( .I1(n22908), .I2(n22907), .O(PE_N18) );
  NR2 U24521 ( .I1(n22910), .I2(n22909), .O(PE_N16) );
  OR2S U24522 ( .I1(n22912), .I2(n22911), .O(n22914) );
  AN2S U24523 ( .I1(n22914), .I2(n22913), .O(PE_N17) );
  INV1S U24524 ( .I(template_store[71]), .O(n23047) );
  INV1S U24525 ( .I(n22915), .O(n22917) );
  NR2 U24526 ( .I1(n23047), .I2(n13914), .O(n22924) );
  NR2 U24527 ( .I1(n23047), .I2(n13915), .O(n23075) );
  INV1S U24528 ( .I(template_store[70]), .O(n23044) );
  NR2 U24529 ( .I1(n23044), .I2(n13914), .O(n23074) );
  NR2 U24530 ( .I1(n23044), .I2(n13915), .O(n23081) );
  NR2 U24531 ( .I1(n23047), .I2(n13916), .O(n23080) );
  INV1S U24532 ( .I(template_store[69]), .O(n23046) );
  NR2 U24533 ( .I1(n23046), .I2(n13914), .O(n23079) );
  OR2S U24534 ( .I1(n22924), .I2(n22925), .O(n23176) );
  ND2S U24535 ( .I1(n22925), .I2(n22924), .O(n23174) );
  ND2S U24536 ( .I1(n23176), .I2(n23174), .O(n23103) );
  INV3 U24537 ( .I(n22929), .O(n23000) );
  NR2 U24538 ( .I1(n23047), .I2(n23000), .O(n22958) );
  NR2 U24539 ( .I1(n23046), .I2(n13912), .O(n22957) );
  INV1S U24540 ( .I(template_store[65]), .O(n23001) );
  NR2 U24541 ( .I1(n23001), .I2(n13915), .O(n22967) );
  INV1S U24542 ( .I(template_store[64]), .O(n23169) );
  NR2 U24543 ( .I1(n23169), .I2(n13914), .O(n22966) );
  INV1S U24544 ( .I(n22933), .O(n22935) );
  NR2 U24545 ( .I1(n23046), .I2(n22936), .O(n22965) );
  INV1S U24546 ( .I(template_store[67]), .O(n23045) );
  NR2 U24547 ( .I1(n23045), .I2(n13916), .O(n22961) );
  INV1S U24548 ( .I(template_store[68]), .O(n23048) );
  INV1S U24549 ( .I(n22937), .O(n22939) );
  NR2 U24550 ( .I1(n23048), .I2(n13925), .O(n22960) );
  NR2 U24551 ( .I1(n23001), .I2(n13914), .O(n22959) );
  INV1S U24552 ( .I(template_store[66]), .O(n22981) );
  NR2 U24553 ( .I1(n22981), .I2(n13916), .O(n22947) );
  NR2 U24554 ( .I1(n23045), .I2(n13925), .O(n22946) );
  NR2 U24555 ( .I1(n23046), .I2(n23000), .O(n22969) );
  NR2 U24556 ( .I1(n23045), .I2(n13912), .O(n22968) );
  NR2 U24557 ( .I1(n22981), .I2(n13915), .O(n22964) );
  NR2 U24558 ( .I1(n23044), .I2(n22936), .O(n22963) );
  NR2 U24559 ( .I1(n23044), .I2(n23000), .O(n22944) );
  NR2 U24560 ( .I1(n23048), .I2(n13912), .O(n22943) );
  NR2 U24561 ( .I1(n23047), .I2(n13913), .O(n22950) );
  HA1 U24562 ( .A(n22944), .B(n22943), .C(n22962), .S(n22949) );
  NR2 U24563 ( .I1(n23001), .I2(n13916), .O(n23017) );
  NR2 U24564 ( .I1(n23044), .I2(n13913), .O(n23016) );
  NR2 U24565 ( .I1(n22981), .I2(n13925), .O(n23015) );
  NR2 U24566 ( .I1(n23169), .I2(n13915), .O(n22972) );
  NR2 U24567 ( .I1(n23048), .I2(n22936), .O(n22971) );
  NR2 U24568 ( .I1(n23048), .I2(n23000), .O(n22986) );
  NR2 U24569 ( .I1(n22981), .I2(n13912), .O(n22985) );
  FA1S U24570 ( .A(n22947), .B(n22946), .CI(n22945), .CO(n22956), .S(n22974)
         );
  FA1S U24571 ( .A(n22950), .B(n22949), .CI(n22948), .CO(n22954), .S(n22973)
         );
  FA1S U24572 ( .A(n22953), .B(n22952), .CI(n22951), .CO(n23069), .S(n22978)
         );
  FA1S U24573 ( .A(n22956), .B(n22955), .CI(n22954), .CO(n23068), .S(n22977)
         );
  NR2 U24574 ( .I1(n23045), .I2(n13915), .O(n23043) );
  NR2 U24575 ( .I1(n22981), .I2(n13914), .O(n23042) );
  NR2 U24576 ( .I1(n23046), .I2(n13925), .O(n23041) );
  NR2 U24577 ( .I1(n23048), .I2(n13916), .O(n23051) );
  NR2 U24578 ( .I1(n23047), .I2(n22936), .O(n23050) );
  HA1 U24579 ( .A(n22958), .B(n22957), .C(n23049), .S(n22953) );
  NR2 U24580 ( .I1(n23044), .I2(n13912), .O(n23060) );
  FA1S U24581 ( .A(n22961), .B(n22960), .CI(n22959), .CO(n23059), .S(n22951)
         );
  FA1S U24582 ( .A(n22964), .B(n22963), .CI(n22962), .CO(n23058), .S(n22955)
         );
  NR2 U24583 ( .I1(n23037), .I2(n23038), .O(n23131) );
  FA1S U24584 ( .A(n22967), .B(n22966), .CI(n22965), .CO(n22952), .S(n23032)
         );
  HA1 U24585 ( .A(n22969), .B(n22968), .C(n22945), .S(n23014) );
  NR2 U24586 ( .I1(n23169), .I2(n13916), .O(n22984) );
  NR2 U24587 ( .I1(n23045), .I2(n22936), .O(n22983) );
  NR2 U24588 ( .I1(n23048), .I2(n13913), .O(n22980) );
  NR2 U24589 ( .I1(n23001), .I2(n13912), .O(n22979) );
  FA1S U24590 ( .A(n22972), .B(n22971), .CI(n22970), .CO(n22975), .S(n23012)
         );
  FA1S U24591 ( .A(n22975), .B(n22974), .CI(n22973), .CO(n22976), .S(n23030)
         );
  FA1S U24592 ( .A(n22978), .B(n22977), .CI(n22976), .CO(n23037), .S(n23036)
         );
  NR2 U24593 ( .I1(n23035), .I2(n23036), .O(n23137) );
  NR2 U24594 ( .I1(n23131), .I2(n23137), .O(n23040) );
  NR2 U24595 ( .I1(n23169), .I2(n13925), .O(n22992) );
  HA1 U24596 ( .A(n22980), .B(n22979), .C(n22982), .S(n22991) );
  NR2 U24597 ( .I1(n23169), .I2(n13912), .O(n22997) );
  NR2 U24598 ( .I1(n23001), .I2(n22936), .O(n22996) );
  NR2 U24599 ( .I1(n22981), .I2(n13913), .O(n22999) );
  NR2 U24600 ( .I1(n23001), .I2(n23000), .O(n22998) );
  NR2 U24601 ( .I1(n23045), .I2(n23000), .O(n22989) );
  NR2 U24602 ( .I1(n22981), .I2(n22936), .O(n22988) );
  NR2 U24603 ( .I1(n22981), .I2(n23000), .O(n22994) );
  NR2 U24604 ( .I1(n23045), .I2(n13913), .O(n22993) );
  FA1S U24605 ( .A(n22984), .B(n22983), .CI(n22982), .CO(n23013), .S(n23022)
         );
  NR2 U24606 ( .I1(n23046), .I2(n13913), .O(n23020) );
  NR2 U24607 ( .I1(n23001), .I2(n13925), .O(n23019) );
  HA1 U24608 ( .A(n22986), .B(n22985), .C(n22970), .S(n23018) );
  NR2 U24609 ( .I1(n23010), .I2(n23011), .O(n23151) );
  FA1S U24610 ( .A(n22989), .B(n22988), .CI(n22987), .CO(n23023), .S(n23007)
         );
  FA1S U24611 ( .A(n22992), .B(n22991), .CI(n22990), .CO(n23010), .S(n23008)
         );
  OR2 U24612 ( .I1(n23007), .I2(n23008), .O(n23157) );
  FA1S U24613 ( .A(n22997), .B(n22996), .CI(n22995), .CO(n22990), .S(n23006)
         );
  NR2 U24614 ( .I1(n23005), .I2(n23006), .O(n23160) );
  NR2 U24615 ( .I1(n23169), .I2(n22936), .O(n23002) );
  HA1 U24616 ( .A(n22999), .B(n22998), .C(n22995), .S(n23003) );
  NR2 U24617 ( .I1(n23169), .I2(n23000), .O(n23170) );
  NR2 U24618 ( .I1(n23001), .I2(n13913), .O(n23171) );
  ND2S U24619 ( .I1(n23170), .I2(n23171), .O(n23172) );
  INV1S U24620 ( .I(n23172), .O(n23168) );
  ND2S U24621 ( .I1(n23003), .I2(n23002), .O(n23165) );
  INV1S U24622 ( .I(n23165), .O(n23004) );
  AOI12HS U24623 ( .B1(n23166), .B2(n23168), .A1(n23004), .O(n23164) );
  OAI12HS U24624 ( .B1(n23160), .B2(n23164), .A1(n23161), .O(n23159) );
  INV1S U24625 ( .I(n23156), .O(n23009) );
  AOI12HS U24626 ( .B1(n23157), .B2(n23159), .A1(n23009), .O(n23155) );
  OAI12HS U24627 ( .B1(n23151), .B2(n23155), .A1(n23152), .O(n23150) );
  FA1S U24628 ( .A(n23014), .B(n23013), .CI(n23012), .CO(n23031), .S(n23024)
         );
  FA1S U24629 ( .A(n23017), .B(n23016), .CI(n23015), .CO(n22948), .S(n23029)
         );
  FA1S U24630 ( .A(n23020), .B(n23019), .CI(n23018), .CO(n23028), .S(n23021)
         );
  FA1S U24631 ( .A(n23023), .B(n23022), .CI(n23021), .CO(n23027), .S(n23011)
         );
  OR2 U24632 ( .I1(n23024), .I2(n23025), .O(n23148) );
  INV1S U24633 ( .I(n23147), .O(n23026) );
  AOI12HS U24634 ( .B1(n23150), .B2(n23148), .A1(n23026), .O(n23146) );
  FA1S U24635 ( .A(n23029), .B(n23028), .CI(n23027), .CO(n23033), .S(n23025)
         );
  FA1S U24636 ( .A(n23032), .B(n23031), .CI(n23030), .CO(n23035), .S(n23034)
         );
  NR2 U24637 ( .I1(n23033), .I2(n23034), .O(n23142) );
  OAI12HS U24638 ( .B1(n23146), .B2(n23142), .A1(n23143), .O(n23134) );
  ND2 U24639 ( .I1(n23036), .I2(n23035), .O(n23138) );
  OAI12HS U24640 ( .B1(n23138), .B2(n23131), .A1(n23132), .O(n23039) );
  AOI12H U24641 ( .B1(n23040), .B2(n23134), .A1(n23039), .O(n23122) );
  NR2 U24642 ( .I1(n23048), .I2(n13915), .O(n23057) );
  NR2 U24643 ( .I1(n23047), .I2(n13912), .O(n23056) );
  FA1S U24644 ( .A(n23043), .B(n23042), .CI(n23041), .CO(n23055), .S(n23066)
         );
  NR2 U24645 ( .I1(n23044), .I2(n13916), .O(n23084) );
  NR2 U24646 ( .I1(n23046), .I2(n13916), .O(n23054) );
  NR2 U24647 ( .I1(n23044), .I2(n13925), .O(n23053) );
  NR2 U24648 ( .I1(n23045), .I2(n13914), .O(n23052) );
  NR2 U24649 ( .I1(n23046), .I2(n13915), .O(n23078) );
  NR2 U24650 ( .I1(n23047), .I2(n13925), .O(n23077) );
  NR2 U24651 ( .I1(n23048), .I2(n13914), .O(n23076) );
  FA1S U24652 ( .A(n23051), .B(n23050), .CI(n23049), .CO(n23063), .S(n23065)
         );
  FA1S U24653 ( .A(n23054), .B(n23053), .CI(n23052), .CO(n23083), .S(n23062)
         );
  FA1S U24654 ( .A(n23057), .B(n23056), .CI(n23055), .CO(n23090), .S(n23061)
         );
  FA1S U24655 ( .A(n23060), .B(n23059), .CI(n23058), .CO(n23072), .S(n23064)
         );
  FA1S U24656 ( .A(n23063), .B(n23062), .CI(n23061), .CO(n23088), .S(n23071)
         );
  FA1S U24657 ( .A(n23066), .B(n23065), .CI(n23064), .CO(n23070), .S(n23067)
         );
  NR2 U24658 ( .I1(n23093), .I2(n23094), .O(n23119) );
  FA1S U24659 ( .A(n23069), .B(n23068), .CI(n23067), .CO(n23091), .S(n23038)
         );
  FA1S U24660 ( .A(n23072), .B(n23071), .CI(n23070), .CO(n23094), .S(n23092)
         );
  NR2 U24661 ( .I1(n23091), .I2(n23092), .O(n23123) );
  NR2 U24662 ( .I1(n23119), .I2(n23123), .O(n23107) );
  FA1S U24663 ( .A(n23075), .B(n23074), .CI(n23073), .CO(n22925), .S(n23097)
         );
  FA1S U24664 ( .A(n23078), .B(n23077), .CI(n23076), .CO(n23087), .S(n23082)
         );
  FA1S U24665 ( .A(n23081), .B(n23080), .CI(n23079), .CO(n23073), .S(n23086)
         );
  FA1S U24666 ( .A(n23084), .B(n23083), .CI(n23082), .CO(n23085), .S(n23089)
         );
  NR2 U24667 ( .I1(n23097), .I2(n23098), .O(n23104) );
  FA1S U24668 ( .A(n23087), .B(n23086), .CI(n23085), .CO(n23098), .S(n23095)
         );
  FA1S U24669 ( .A(n23090), .B(n23089), .CI(n23088), .CO(n23096), .S(n23093)
         );
  NR2 U24670 ( .I1(n23095), .I2(n23096), .O(n23111) );
  NR2 U24671 ( .I1(n23104), .I2(n23111), .O(n23100) );
  ND2 U24672 ( .I1(n23092), .I2(n23091), .O(n23127) );
  OAI12HS U24673 ( .B1(n23119), .B2(n23127), .A1(n23120), .O(n23108) );
  OAI12HS U24674 ( .B1(n23115), .B2(n23104), .A1(n23105), .O(n23099) );
  AOI12HS U24675 ( .B1(n23108), .B2(n23100), .A1(n23099), .O(n23101) );
  OAI12HS U24676 ( .B1(n23122), .B2(n23102), .A1(n23101), .O(n23177) );
  XNR2HS U24677 ( .I1(n23103), .I2(n23177), .O(PE_N14) );
  INV1S U24678 ( .I(n23104), .O(n23106) );
  ND2S U24679 ( .I1(n23106), .I2(n23105), .O(n23114) );
  INV1S U24680 ( .I(n23107), .O(n23110) );
  INV1S U24681 ( .I(n23108), .O(n23109) );
  INV1S U24682 ( .I(n23111), .O(n23116) );
  INV1S U24683 ( .I(n23115), .O(n23112) );
  AOI12HS U24684 ( .B1(n23117), .B2(n23116), .A1(n23112), .O(n23113) );
  XOR2HS U24685 ( .I1(n23114), .I2(n23113), .O(PE_N13) );
  ND2S U24686 ( .I1(n23116), .I2(n23115), .O(n23118) );
  XNR2HS U24687 ( .I1(n23118), .I2(n23117), .O(PE_N12) );
  INV1S U24688 ( .I(n23119), .O(n23121) );
  INV1S U24689 ( .I(n23123), .O(n23128) );
  INV1S U24690 ( .I(n23127), .O(n23124) );
  AOI12HS U24691 ( .B1(n23129), .B2(n23128), .A1(n23124), .O(n23125) );
  XOR2HS U24692 ( .I1(n23126), .I2(n23125), .O(PE_N11) );
  XNR2HS U24693 ( .I1(n23130), .I2(n23129), .O(PE_N10) );
  INV1S U24694 ( .I(n23131), .O(n23133) );
  INV1S U24695 ( .I(n23134), .O(n23141) );
  OAI12HS U24696 ( .B1(n23141), .B2(n23137), .A1(n23138), .O(n23135) );
  XNR2HS U24697 ( .I1(n23136), .I2(n23135), .O(PE_N9) );
  INV1S U24698 ( .I(n23137), .O(n23139) );
  XOR2HS U24699 ( .I1(n23141), .I2(n23140), .O(PE_N8) );
  INV1S U24700 ( .I(n23142), .O(n23144) );
  ND2S U24701 ( .I1(n23144), .I2(n23143), .O(n23145) );
  XOR2HS U24702 ( .I1(n23146), .I2(n23145), .O(PE_N7) );
  ND2S U24703 ( .I1(n23148), .I2(n23147), .O(n23149) );
  XNR2HS U24704 ( .I1(n23150), .I2(n23149), .O(PE_N6) );
  INV1S U24705 ( .I(n23151), .O(n23153) );
  ND2S U24706 ( .I1(n23153), .I2(n23152), .O(n23154) );
  XOR2HS U24707 ( .I1(n23155), .I2(n23154), .O(PE_N5) );
  ND2S U24708 ( .I1(n23157), .I2(n23156), .O(n23158) );
  XNR2HS U24709 ( .I1(n23159), .I2(n23158), .O(PE_N4) );
  INV1S U24710 ( .I(n23160), .O(n23162) );
  ND2S U24711 ( .I1(n23162), .I2(n23161), .O(n23163) );
  XOR2HS U24712 ( .I1(n23164), .I2(n23163), .O(PE_N3) );
  ND2S U24713 ( .I1(n23166), .I2(n23165), .O(n23167) );
  XNR2HS U24714 ( .I1(n23168), .I2(n23167), .O(PE_N2) );
  NR2 U24715 ( .I1(n23169), .I2(n13913), .O(PE_N0) );
  OR2S U24716 ( .I1(n23171), .I2(n23170), .O(n23173) );
  AN2S U24717 ( .I1(n23173), .I2(n23172), .O(PE_N1) );
  INV1S U24718 ( .I(n23174), .O(n23175) );
  AO12 U24719 ( .B1(n23177), .B2(n23176), .A1(n23175), .O(PE_N15) );
  INV1S U24720 ( .I(template_store[55]), .O(n23300) );
  NR2 U24721 ( .I1(n23300), .I2(n23292), .O(n23181) );
  INV1S U24722 ( .I(template_store[54]), .O(n23296) );
  NR2 U24723 ( .I1(n23296), .I2(n23292), .O(n23345) );
  NR2 U24724 ( .I1(n23300), .I2(n23297), .O(n23344) );
  NR2 U24725 ( .I1(n23300), .I2(n23295), .O(n23336) );
  INV1S U24726 ( .I(template_store[53]), .O(n23298) );
  NR2 U24727 ( .I1(n23298), .I2(n23292), .O(n23335) );
  NR2 U24728 ( .I1(n23296), .I2(n23297), .O(n23334) );
  NR2 U24729 ( .I1(n23181), .I2(n23182), .O(n23361) );
  INV1S U24730 ( .I(n23361), .O(n23183) );
  ND2S U24731 ( .I1(n23182), .I2(n23181), .O(n23360) );
  ND2S U24732 ( .I1(n23183), .I2(n23360), .O(n23357) );
  INV1S U24733 ( .I(template_store[50]), .O(n23225) );
  NR2 U24734 ( .I1(n23225), .I2(n23299), .O(n23191) );
  INV1S U24735 ( .I(template_store[51]), .O(n23288) );
  NR2 U24736 ( .I1(n23288), .I2(n23294), .O(n23190) );
  INV1S U24737 ( .I(template_store[49]), .O(n23248) );
  NR2 U24738 ( .I1(n23248), .I2(n23295), .O(n23193) );
  INV1S U24739 ( .I(template_store[48]), .O(n23428) );
  NR2 U24740 ( .I1(n23428), .I2(n23297), .O(n23192) );
  INV1S U24741 ( .I(template_store[52]), .O(n23293) );
  NR2 U24742 ( .I1(n23293), .I2(n23244), .O(n23261) );
  INV2 U24743 ( .I(n23187), .O(n23427) );
  NR2 U24744 ( .I1(n23298), .I2(n23427), .O(n23230) );
  NR2 U24745 ( .I1(n23288), .I2(n23244), .O(n23229) );
  NR2 U24746 ( .I1(n23428), .I2(n23299), .O(n23232) );
  INV2 U24747 ( .I(n23188), .O(n23247) );
  NR2 U24748 ( .I1(n23288), .I2(n23247), .O(n23231) );
  FA1S U24749 ( .A(n23191), .B(n23190), .CI(n23189), .CO(n23279), .S(n23259)
         );
  NR2 U24750 ( .I1(n23248), .I2(n23297), .O(n23202) );
  NR2 U24751 ( .I1(n23300), .I2(n23427), .O(n23201) );
  NR2 U24752 ( .I1(n23225), .I2(n23295), .O(n23204) );
  NR2 U24753 ( .I1(n23428), .I2(n23292), .O(n23203) );
  NR2 U24754 ( .I1(n23288), .I2(n23299), .O(n23196) );
  NR2 U24755 ( .I1(n23293), .I2(n23294), .O(n23195) );
  NR2 U24756 ( .I1(n23296), .I2(n23247), .O(n23207) );
  NR2 U24757 ( .I1(n23298), .I2(n23244), .O(n23206) );
  NR2 U24758 ( .I1(n23298), .I2(n23247), .O(n23264) );
  NR2 U24759 ( .I1(n23296), .I2(n23427), .O(n23263) );
  NR2 U24760 ( .I1(n23428), .I2(n23295), .O(n23227) );
  NR2 U24761 ( .I1(n23248), .I2(n23299), .O(n23226) );
  NR2 U24762 ( .I1(n23296), .I2(n23244), .O(n23224) );
  FA1S U24763 ( .A(n23196), .B(n23195), .CI(n23194), .CO(n23223), .S(n23198)
         );
  NR2 U24764 ( .I1(n23225), .I2(n23297), .O(n23221) );
  NR2 U24765 ( .I1(n23300), .I2(n23247), .O(n23220) );
  NR2 U24766 ( .I1(n23288), .I2(n23295), .O(n23215) );
  NR2 U24767 ( .I1(n23248), .I2(n23292), .O(n23214) );
  FA1S U24768 ( .A(n23199), .B(n23198), .CI(n23197), .CO(n23209), .S(n23277)
         );
  FA1S U24769 ( .A(n23202), .B(n23201), .CI(n23200), .CO(n23218), .S(n23199)
         );
  NR2 U24770 ( .I1(n23293), .I2(n23299), .O(n23213) );
  NR2 U24771 ( .I1(n23298), .I2(n23294), .O(n23212) );
  FA1S U24772 ( .A(n23207), .B(n23206), .CI(n23205), .CO(n23216), .S(n23197)
         );
  NR2 U24773 ( .I1(n23282), .I2(n23283), .O(n23395) );
  FA1S U24774 ( .A(n23210), .B(n23209), .CI(n23208), .CO(n23284), .S(n23283)
         );
  NR2 U24775 ( .I1(n23296), .I2(n23294), .O(n23312) );
  FA1S U24776 ( .A(n23213), .B(n23212), .CI(n23211), .CO(n23311), .S(n23217)
         );
  NR2 U24777 ( .I1(n23293), .I2(n23295), .O(n23303) );
  NR2 U24778 ( .I1(n23298), .I2(n23299), .O(n23302) );
  FA1S U24779 ( .A(n23218), .B(n23217), .CI(n23216), .CO(n23320), .S(n23208)
         );
  NR2 U24780 ( .I1(n23225), .I2(n23292), .O(n23291) );
  NR2 U24781 ( .I1(n23288), .I2(n23297), .O(n23290) );
  NR2 U24782 ( .I1(n23300), .I2(n23244), .O(n23289) );
  FA1S U24783 ( .A(n23221), .B(n23220), .CI(n23219), .CO(n23317), .S(n23222)
         );
  FA1S U24784 ( .A(n23224), .B(n23223), .CI(n23222), .CO(n23316), .S(n23210)
         );
  NR2 U24785 ( .I1(n23395), .I2(n23389), .O(n23287) );
  NR2 U24786 ( .I1(n23225), .I2(n23244), .O(n23238) );
  NR2 U24787 ( .I1(n23288), .I2(n23427), .O(n23240) );
  NR2 U24788 ( .I1(n23225), .I2(n23247), .O(n23239) );
  NR2 U24789 ( .I1(n23428), .I2(n23294), .O(n23243) );
  NR2 U24790 ( .I1(n23248), .I2(n23244), .O(n23242) );
  NR2 U24791 ( .I1(n23225), .I2(n23427), .O(n23246) );
  NR2 U24792 ( .I1(n23248), .I2(n23247), .O(n23245) );
  NR2 U24793 ( .I1(n23293), .I2(n23247), .O(n23267) );
  NR2 U24794 ( .I1(n23225), .I2(n23294), .O(n23266) );
  HA1 U24795 ( .A(n23227), .B(n23226), .C(n23262), .S(n23265) );
  FA1S U24796 ( .A(n23230), .B(n23229), .CI(n23228), .CO(n23260), .S(n23269)
         );
  NR2 U24797 ( .I1(n23293), .I2(n23427), .O(n23235) );
  NR2 U24798 ( .I1(n23248), .I2(n23294), .O(n23234) );
  NR2 U24799 ( .I1(n23257), .I2(n23258), .O(n23409) );
  FA1S U24800 ( .A(n23235), .B(n23234), .CI(n23233), .CO(n23268), .S(n23254)
         );
  FA1S U24801 ( .A(n23238), .B(n23237), .CI(n23236), .CO(n23257), .S(n23255)
         );
  OR2 U24802 ( .I1(n23254), .I2(n23255), .O(n23415) );
  FA1S U24803 ( .A(n23243), .B(n23242), .CI(n23241), .CO(n23236), .S(n23253)
         );
  NR2 U24804 ( .I1(n23252), .I2(n23253), .O(n23418) );
  NR2 U24805 ( .I1(n23428), .I2(n23244), .O(n23249) );
  NR2 U24806 ( .I1(n23428), .I2(n23247), .O(n23429) );
  NR2 U24807 ( .I1(n23248), .I2(n23427), .O(n23430) );
  ND2S U24808 ( .I1(n23429), .I2(n23430), .O(n23431) );
  INV1S U24809 ( .I(n23431), .O(n23426) );
  ND2S U24810 ( .I1(n23250), .I2(n23249), .O(n23423) );
  INV1S U24811 ( .I(n23423), .O(n23251) );
  AOI12HS U24812 ( .B1(n23424), .B2(n23426), .A1(n23251), .O(n23422) );
  ND2S U24813 ( .I1(n23253), .I2(n23252), .O(n23419) );
  OAI12HS U24814 ( .B1(n23418), .B2(n23422), .A1(n23419), .O(n23417) );
  INV1S U24815 ( .I(n23414), .O(n23256) );
  AOI12HS U24816 ( .B1(n23415), .B2(n23417), .A1(n23256), .O(n23413) );
  OAI12HS U24817 ( .B1(n23409), .B2(n23413), .A1(n23410), .O(n23407) );
  FA1S U24818 ( .A(n23261), .B(n23260), .CI(n23259), .CO(n23278), .S(n23271)
         );
  FA1S U24819 ( .A(n23264), .B(n23263), .CI(n23262), .CO(n23205), .S(n23276)
         );
  FA1S U24820 ( .A(n23267), .B(n23266), .CI(n23265), .CO(n23275), .S(n23270)
         );
  FA1S U24821 ( .A(n23270), .B(n23269), .CI(n23268), .CO(n23274), .S(n23258)
         );
  OR2 U24822 ( .I1(n23271), .I2(n23272), .O(n23406) );
  INV1S U24823 ( .I(n23405), .O(n23273) );
  AOI12HS U24824 ( .B1(n23407), .B2(n23406), .A1(n23273), .O(n23403) );
  FA1S U24825 ( .A(n23276), .B(n23275), .CI(n23274), .CO(n23280), .S(n23272)
         );
  FA1S U24826 ( .A(n23279), .B(n23278), .CI(n23277), .CO(n23282), .S(n23281)
         );
  NR2 U24827 ( .I1(n23280), .I2(n23281), .O(n23400) );
  OAI12HS U24828 ( .B1(n23403), .B2(n23400), .A1(n23401), .O(n23392) );
  ND2 U24829 ( .I1(n23283), .I2(n23282), .O(n23396) );
  ND2 U24830 ( .I1(n23285), .I2(n23284), .O(n23390) );
  OAI12HS U24831 ( .B1(n23389), .B2(n23396), .A1(n23390), .O(n23286) );
  AOI12H U24832 ( .B1(n23287), .B2(n23392), .A1(n23286), .O(n23380) );
  NR2 U24833 ( .I1(n23288), .I2(n23292), .O(n23309) );
  NR2 U24834 ( .I1(n23293), .I2(n23297), .O(n23308) );
  FA1S U24835 ( .A(n23291), .B(n23290), .CI(n23289), .CO(n23307), .S(n23318)
         );
  NR2 U24836 ( .I1(n23293), .I2(n23292), .O(n23339) );
  NR2 U24837 ( .I1(n23298), .I2(n23295), .O(n23306) );
  NR2 U24838 ( .I1(n23296), .I2(n23299), .O(n23305) );
  NR2 U24839 ( .I1(n23300), .I2(n23294), .O(n23304) );
  NR2 U24840 ( .I1(n23296), .I2(n23295), .O(n23333) );
  NR2 U24841 ( .I1(n23298), .I2(n23297), .O(n23332) );
  NR2 U24842 ( .I1(n23300), .I2(n23299), .O(n23331) );
  FA1S U24843 ( .A(n23303), .B(n23302), .CI(n23301), .CO(n23315), .S(n23310)
         );
  FA1S U24844 ( .A(n23306), .B(n23305), .CI(n23304), .CO(n23338), .S(n23314)
         );
  FA1S U24845 ( .A(n23309), .B(n23308), .CI(n23307), .CO(n23342), .S(n23313)
         );
  FA1S U24846 ( .A(n23312), .B(n23311), .CI(n23310), .CO(n23324), .S(n23321)
         );
  FA1S U24847 ( .A(n23315), .B(n23314), .CI(n23313), .CO(n23340), .S(n23323)
         );
  FA1S U24848 ( .A(n23318), .B(n23317), .CI(n23316), .CO(n23322), .S(n23319)
         );
  NR2 U24849 ( .I1(n23327), .I2(n23328), .O(n23377) );
  FA1 U24850 ( .A(n23321), .B(n23320), .CI(n23319), .CO(n23325), .S(n23285) );
  NR2 U24851 ( .I1(n23325), .I2(n23326), .O(n23381) );
  NR2 U24852 ( .I1(n23377), .I2(n23381), .O(n23359) );
  INV1S U24853 ( .I(n23359), .O(n23330) );
  ND2 U24854 ( .I1(n23328), .I2(n23327), .O(n23378) );
  OAI12HS U24855 ( .B1(n23377), .B2(n23385), .A1(n23378), .O(n23365) );
  INV1S U24856 ( .I(n23365), .O(n23329) );
  FA1S U24857 ( .A(n23333), .B(n23332), .CI(n23331), .CO(n23348), .S(n23337)
         );
  FA1S U24858 ( .A(n23336), .B(n23335), .CI(n23334), .CO(n23343), .S(n23347)
         );
  FA1S U24859 ( .A(n23339), .B(n23338), .CI(n23337), .CO(n23346), .S(n23341)
         );
  FA1S U24860 ( .A(n23342), .B(n23341), .CI(n23340), .CO(n23350), .S(n23327)
         );
  OR2 U24861 ( .I1(n23349), .I2(n23350), .O(n23374) );
  FA1S U24862 ( .A(n23345), .B(n23344), .CI(n23343), .CO(n23182), .S(n23351)
         );
  FA1S U24863 ( .A(n23348), .B(n23347), .CI(n23346), .CO(n23352), .S(n23349)
         );
  INV1S U24864 ( .I(n23358), .O(n23355) );
  INV1S U24865 ( .I(n23373), .O(n23370) );
  INV1S U24866 ( .I(n23368), .O(n23353) );
  AOI12HS U24867 ( .B1(n23370), .B2(n23369), .A1(n23353), .O(n23362) );
  INV1S U24868 ( .I(n23362), .O(n23354) );
  AOI12HS U24869 ( .B1(n23375), .B2(n23355), .A1(n23354), .O(n23356) );
  XOR2HS U24870 ( .I1(n23357), .I2(n23356), .O(PE_N46) );
  NR2 U24871 ( .I1(n23361), .I2(n23358), .O(n23364) );
  OAI12HS U24872 ( .B1(n23362), .B2(n23361), .A1(n23360), .O(n23363) );
  AOI12HS U24873 ( .B1(n23365), .B2(n23364), .A1(n23363), .O(n23366) );
  OAI12HS U24874 ( .B1(n23380), .B2(n23367), .A1(n23366), .O(PE_N47) );
  ND2S U24875 ( .I1(n23369), .I2(n23368), .O(n23372) );
  AOI12HS U24876 ( .B1(n23375), .B2(n23374), .A1(n23370), .O(n23371) );
  XOR2HS U24877 ( .I1(n23372), .I2(n23371), .O(PE_N45) );
  ND2S U24878 ( .I1(n23374), .I2(n23373), .O(n23376) );
  XNR2HS U24879 ( .I1(n23376), .I2(n23375), .O(PE_N44) );
  INV1S U24880 ( .I(n23377), .O(n23379) );
  INV1S U24881 ( .I(n23381), .O(n23386) );
  INV1S U24882 ( .I(n23385), .O(n23382) );
  AOI12HS U24883 ( .B1(n23387), .B2(n23386), .A1(n23382), .O(n23383) );
  XOR2HS U24884 ( .I1(n23384), .I2(n23383), .O(PE_N43) );
  XNR2HS U24885 ( .I1(n23388), .I2(n23387), .O(PE_N42) );
  INV1S U24886 ( .I(n23389), .O(n23391) );
  ND2S U24887 ( .I1(n23391), .I2(n23390), .O(n23394) );
  INV1S U24888 ( .I(n23392), .O(n23399) );
  OAI12HS U24889 ( .B1(n23399), .B2(n23395), .A1(n23396), .O(n23393) );
  XNR2HS U24890 ( .I1(n23394), .I2(n23393), .O(PE_N41) );
  INV1S U24891 ( .I(n23395), .O(n23397) );
  XOR2HS U24892 ( .I1(n23399), .I2(n23398), .O(PE_N40) );
  INV1S U24893 ( .I(n23400), .O(n23402) );
  ND2S U24894 ( .I1(n23402), .I2(n23401), .O(n23404) );
  XOR2HS U24895 ( .I1(n23404), .I2(n23403), .O(PE_N39) );
  ND2S U24896 ( .I1(n23406), .I2(n23405), .O(n23408) );
  XNR2HS U24897 ( .I1(n23408), .I2(n23407), .O(PE_N38) );
  INV1S U24898 ( .I(n23409), .O(n23411) );
  ND2S U24899 ( .I1(n23411), .I2(n23410), .O(n23412) );
  XOR2HS U24900 ( .I1(n23413), .I2(n23412), .O(PE_N37) );
  ND2S U24901 ( .I1(n23415), .I2(n23414), .O(n23416) );
  XNR2HS U24902 ( .I1(n23417), .I2(n23416), .O(PE_N36) );
  INV1S U24903 ( .I(n23418), .O(n23420) );
  ND2S U24904 ( .I1(n23420), .I2(n23419), .O(n23421) );
  XOR2HS U24905 ( .I1(n23422), .I2(n23421), .O(PE_N35) );
  ND2S U24906 ( .I1(n23424), .I2(n23423), .O(n23425) );
  XNR2HS U24907 ( .I1(n23426), .I2(n23425), .O(PE_N34) );
  NR2 U24908 ( .I1(n23428), .I2(n23427), .O(PE_N32) );
  OR2S U24909 ( .I1(n23430), .I2(n23429), .O(n23432) );
  AN2S U24910 ( .I1(n23432), .I2(n23431), .O(PE_N33) );
  INV1S U24911 ( .I(n23433), .O(n23435) );
  ND2S U24912 ( .I1(n23435), .I2(n23434), .O(n23436) );
  XOR2HS U24913 ( .I1(n23437), .I2(n23436), .O(n23455) );
  INV1S U24914 ( .I(n23455), .O(n23454) );
  NR2 U24915 ( .I1(n23454), .I2(n23445), .O(n23439) );
  NR2 U24916 ( .I1(n23439), .I2(n23438), .O(n23443) );
  INV1S U24917 ( .I(n23440), .O(n23441) );
  INV1S U24918 ( .I(gray_avg[3]), .O(n23444) );
  AOI22S U24919 ( .A1(gray_avg[3]), .A2(n23445), .B1(n23444), .B2(n23446), .O(
        n23450) );
  AN2B1S U24920 ( .I1(n23445), .B1(n23454), .O(n23448) );
  XOR2HS U24921 ( .I1(n23454), .I2(n23446), .O(n23447) );
  MXL2HS U24922 ( .A(n23448), .B(n23447), .S(gray_avg[3]), .OB(n23449) );
  MXL2HS U24923 ( .A(n23450), .B(n23449), .S(gray_avg[2]), .OB(n23465) );
  ND2S U24924 ( .I1(n13928), .I2(n23451), .O(n23452) );
  INV1S U24925 ( .I(n23463), .O(n23457) );
  NR2 U24926 ( .I1(n13921), .I2(n23457), .O(n23458) );
  INV1S U24927 ( .I(n23459), .O(n23461) );
  ND2S U24928 ( .I1(n23461), .I2(n23460), .O(n23462) );
  NR2 U24929 ( .I1(n13920), .I2(n13921), .O(n23464) );
  INV1S U24930 ( .I(n23465), .O(n23466) );
  NR2 U24931 ( .I1(n13917), .I2(n23466), .O(n23467) );
  NR2 U24932 ( .I1(n23470), .I2(n22942), .O(PE_N64) );
  NR2 U24933 ( .I1(n23526), .I2(n13817), .O(n23486) );
  NR2 U24934 ( .I1(n23509), .I2(n23508), .O(n23485) );
  FA1S U24935 ( .A(n23473), .B(n23472), .CI(n23471), .CO(n23484), .S(n23476)
         );
  FA1S U24936 ( .A(n23476), .B(n23475), .CI(n23474), .CO(n23498), .S(n23494)
         );
  FA1S U24937 ( .A(n23479), .B(n23478), .CI(n23477), .CO(n23493), .S(n23481)
         );
  NR2 U24938 ( .I1(n23536), .I2(n13816), .O(n23489) );
  NR2 U24939 ( .I1(n23537), .I2(n23480), .O(n23488) );
  NR2 U24940 ( .I1(n23490), .I2(n23525), .O(n23487) );
  FA1S U24941 ( .A(n23483), .B(n23482), .CI(n23481), .CO(n23491), .S(n23496)
         );
  FA1S U24942 ( .A(n23486), .B(n23485), .CI(n23484), .CO(n23515), .S(n23499)
         );
  NR2 U24943 ( .I1(n23526), .I2(n23508), .O(n23512) );
  FA1S U24944 ( .A(n23489), .B(n23488), .CI(n23487), .CO(n23511), .S(n23492)
         );
  NR2 U24945 ( .I1(n23536), .I2(n13817), .O(n23507) );
  NR2 U24946 ( .I1(n23537), .I2(n23490), .O(n23506) );
  NR2 U24947 ( .I1(n23509), .I2(n23525), .O(n23505) );
  FA1S U24948 ( .A(n23493), .B(n23492), .CI(n23491), .CO(n23513), .S(n23497)
         );
  FA1S U24949 ( .A(n23496), .B(n23495), .CI(n23494), .CO(n23521), .S(n23502)
         );
  FA1S U24950 ( .A(n23499), .B(n23498), .CI(n23497), .CO(n23518), .S(n23520)
         );
  INV1S U24951 ( .I(n23500), .O(n23504) );
  FA1S U24952 ( .A(n23507), .B(n23506), .CI(n23505), .CO(n23532), .S(n23510)
         );
  NR2 U24953 ( .I1(n23536), .I2(n23508), .O(n23529) );
  NR2 U24954 ( .I1(n23537), .I2(n23509), .O(n23528) );
  NR2 U24955 ( .I1(n23526), .I2(n23525), .O(n23527) );
  FA1S U24956 ( .A(n23512), .B(n23511), .CI(n23510), .CO(n23530), .S(n23514)
         );
  FA1S U24957 ( .A(n23515), .B(n23514), .CI(n23513), .CO(n23534), .S(n23517)
         );
  FA1 U24958 ( .A(n23518), .B(n23517), .CI(n23516), .CO(n23533), .S(PE_N75) );
  FA1 U24959 ( .A(n23521), .B(n23520), .CI(n23519), .CO(n23516), .S(PE_N74) );
  FA1 U24960 ( .A(n23524), .B(n23523), .CI(n23522), .CO(n23500), .S(PE_N72) );
  NR2 U24961 ( .I1(n23536), .I2(n23525), .O(n23540) );
  NR2 U24962 ( .I1(n23537), .I2(n23526), .O(n23539) );
  FA1S U24963 ( .A(n23529), .B(n23528), .CI(n23527), .CO(n23538), .S(n23531)
         );
  FA1S U24964 ( .A(n23532), .B(n23531), .CI(n23530), .CO(n23542), .S(n23535)
         );
  FA1 U24965 ( .A(n23535), .B(n23534), .CI(n23533), .CO(n23541), .S(PE_N76) );
  NR2 U24966 ( .I1(n23537), .I2(n23536), .O(n23546) );
  FA1S U24967 ( .A(n23540), .B(n23539), .CI(n23538), .CO(n23545), .S(n23543)
         );
  FA1 U24968 ( .A(n23543), .B(n23542), .CI(n23541), .CO(n23544), .S(PE_N77) );
  FA1 U24969 ( .A(n23546), .B(n23545), .CI(n23544), .CO(PE_N79), .S(PE_N78) );
  FA1 U24970 ( .A(n23549), .B(n23548), .CI(n23547), .CO(n23550), .S(PE_N69) );
  FA1 U24971 ( .A(n23552), .B(n23551), .CI(n23550), .CO(n21630), .S(PE_N70) );
  FA1 U24972 ( .A(n23555), .B(n23554), .CI(n23553), .CO(n21724), .S(PE_N66) );
  FA1 U24973 ( .A(n23558), .B(n23557), .CI(n23556), .CO(n23547), .S(PE_N68) );
  OR2T U24974 ( .I1(n23559), .I2(n30028), .O(n23808) );
  NR2P U24975 ( .I1(n23640), .I2(n23808), .O(n30039) );
  INV1S U24976 ( .I(n23808), .O(n30036) );
  BUF1 U24977 ( .I(n13805), .O(n30034) );
  BUF1 U24978 ( .I(rst_n), .O(n30035) );
  INV1S U24979 ( .I(addr[2]), .O(n30007) );
  ND2S U24980 ( .I1(addr[1]), .I2(addr[0]), .O(n30005) );
  NR2 U24981 ( .I1(n30007), .I2(n30005), .O(n30008) );
  ND2S U24982 ( .I1(addr[3]), .I2(n30008), .O(n30012) );
  NR2 U24983 ( .I1(n23560), .I2(n30012), .O(n30018) );
  INV1S U24984 ( .I(in_cnt[1]), .O(n29958) );
  INV1S U24985 ( .I(in_cnt[0]), .O(n29960) );
  ND2S U24986 ( .I1(n29958), .I2(n29960), .O(n23564) );
  OR2S U24987 ( .I1(N25894), .I2(n23564), .O(n23562) );
  ND2S U24988 ( .I1(n23562), .I2(n23561), .O(n30014) );
  ND3S U24989 ( .I1(addr[6]), .I2(n30018), .I3(n30014), .O(n23567) );
  ND2S U24990 ( .I1(addr[6]), .I2(n30018), .O(n23563) );
  ND2S U24991 ( .I1(n30014), .I2(n23563), .O(n23566) );
  AOI13HS U24992 ( .B1(c_s[0]), .B2(n23565), .B3(n23564), .A1(c_s[2]), .O(
        n30011) );
  ND2S U24993 ( .I1(n23566), .I2(n30011), .O(n23616) );
  MOAI1S U24994 ( .A1(addr[7]), .A2(n23567), .B1(addr[7]), .B2(n23616), .O(
        n13633) );
  INV1S U24995 ( .I(rgb_value[11]), .O(n29930) );
  INV1S U24996 ( .I(rgb_value[20]), .O(n29929) );
  ND2S U24997 ( .I1(n29929), .I2(n29930), .O(n23568) );
  MOAI1S U24998 ( .A1(n29930), .A2(n29929), .B1(n23568), .B2(rgb_value[4]), 
        .O(intadd_8_A_3_) );
  INV1S U24999 ( .I(rgb_value[12]), .O(n29928) );
  INV1S U25000 ( .I(rgb_value[21]), .O(n29927) );
  ND2S U25001 ( .I1(n29927), .I2(n29928), .O(n23569) );
  MOAI1S U25002 ( .A1(n29928), .A2(n29927), .B1(n23569), .B2(rgb_value[5]), 
        .O(intadd_8_B_4_) );
  INV1S U25003 ( .I(rgb_value[13]), .O(n29926) );
  INV1S U25004 ( .I(rgb_value[22]), .O(n29925) );
  ND2S U25005 ( .I1(n29925), .I2(n29926), .O(n23570) );
  MOAI1S U25006 ( .A1(n29926), .A2(n29925), .B1(n23570), .B2(rgb_value[6]), 
        .O(intadd_8_B_5_) );
  NR2 U25007 ( .I1(n23572), .I2(n23571), .O(n23573) );
  ND2S U25008 ( .I1(n23573), .I2(image_size[0]), .O(n23664) );
  INV1S U25009 ( .I(n23573), .O(n23666) );
  MOAI1S U25010 ( .A1(image_size[1]), .A2(n23664), .B1(n23666), .B2(
        img_size_hold[3]), .O(n11202) );
  INV1S U25011 ( .I(action[2]), .O(n23575) );
  INV1S U25012 ( .I(act_cnt[0]), .O(n29966) );
  NR2 U25013 ( .I1(n29962), .I2(n29966), .O(n23651) );
  INV1S U25014 ( .I(act_cnt[2]), .O(n23649) );
  INV1S U25015 ( .I(act_cnt[1]), .O(n29964) );
  INV1S U25016 ( .I(n23652), .O(n23581) );
  INV1S U25017 ( .I(n23578), .O(n23574) );
  NR2 U25018 ( .I1(n23581), .I2(n23574), .O(n23577) );
  MOAI1S U25019 ( .A1(n23575), .A2(n23578), .B1(n23577), .B2(act[20]), .O(
        n13659) );
  INV1S U25020 ( .I(action[0]), .O(n23576) );
  MOAI1S U25021 ( .A1(n23576), .A2(n23578), .B1(n23577), .B2(act[18]), .O(
        n13660) );
  INV1S U25022 ( .I(action[1]), .O(n23579) );
  MOAI1S U25023 ( .A1(n23579), .A2(n23578), .B1(n23577), .B2(act[19]), .O(
        n13658) );
  INV1S U25024 ( .I(n23655), .O(n23582) );
  ND3S U25025 ( .I1(n23651), .I2(act_cnt[1]), .I3(n23649), .O(n23628) );
  INV1S U25026 ( .I(n23628), .O(n23580) );
  NR2 U25027 ( .I1(n23581), .I2(n23580), .O(n23584) );
  MOAI1S U25028 ( .A1(n23582), .A2(n23628), .B1(n23584), .B2(act[14]), .O(
        n13665) );
  INV1S U25029 ( .I(n23654), .O(n23583) );
  MOAI1S U25030 ( .A1(n23583), .A2(n23628), .B1(n23584), .B2(act[13]), .O(
        n13664) );
  INV1S U25031 ( .I(n23663), .O(n23585) );
  MOAI1S U25032 ( .A1(n23585), .A2(n23628), .B1(n23584), .B2(act[12]), .O(
        n13666) );
  INV1S U25033 ( .I(n23682), .O(n23675) );
  NR2 U25034 ( .I1(n29996), .I2(n29999), .O(n29995) );
  AN3B2S U25035 ( .I1(n23587), .B1(n23586), .B2(n30029), .O(n30021) );
  INV1S U25036 ( .I(n30021), .O(n29998) );
  OA112S U25037 ( .C1(set_cnt[1]), .C2(n29995), .A1(n29997), .B1(n29998), .O(
        n13636) );
  NR2 U25038 ( .I1(n23900), .I2(img_size[1]), .O(n23591) );
  ND2S U25039 ( .I1(n23591), .I2(n23932), .O(n23698) );
  OR2S U25040 ( .I1(n23932), .I2(n23591), .O(n23588) );
  AN2S U25041 ( .I1(n23698), .I2(n23588), .O(n23749) );
  OR2S U25042 ( .I1(i_col[3]), .I2(n23749), .O(n23590) );
  XNR2HS U25043 ( .I1(n23589), .I2(n23698), .O(n23751) );
  ND3S U25044 ( .I1(n23590), .I2(n23665), .I3(n23751), .O(n23804) );
  INV1S U25045 ( .I(n23804), .O(n23596) );
  INV1S U25046 ( .I(n23860), .O(n23922) );
  NR2 U25047 ( .I1(n23591), .I2(n23922), .O(n23701) );
  ND2S U25048 ( .I1(n23701), .I2(i_col[2]), .O(n23805) );
  OR2S U25049 ( .I1(i_col[2]), .I2(n23701), .O(n23803) );
  ND2S U25050 ( .I1(i_col[1]), .I2(img_size[1]), .O(n23800) );
  OAI12HS U25051 ( .B1(n28555), .B2(n23592), .A1(n23800), .O(n23593) );
  OAI22S U25052 ( .A1(i_col[0]), .A2(n28540), .B1(i_col[1]), .B2(img_size[1]), 
        .O(n23801) );
  NR2 U25053 ( .I1(n23593), .I2(n23801), .O(n23594) );
  AN3S U25054 ( .I1(n23805), .I2(n23803), .I3(n23594), .O(n23595) );
  ND2S U25055 ( .I1(n23749), .I2(i_col[3]), .O(n23807) );
  ND3S U25056 ( .I1(n23596), .I2(n23595), .I3(n23807), .O(n23598) );
  NR2 U25057 ( .I1(n29968), .I2(n23607), .O(n23812) );
  NR2 U25058 ( .I1(n24698), .I2(n23698), .O(n24043) );
  INV1S U25059 ( .I(n24043), .O(n23597) );
  ND2S U25060 ( .I1(n23812), .I2(n23597), .O(n23699) );
  NR2 U25061 ( .I1(n23598), .I2(n23699), .O(n23603) );
  INV1S U25062 ( .I(n23603), .O(n23622) );
  NR2 U25063 ( .I1(n23827), .I2(n23622), .O(n23830) );
  NR3 U25064 ( .I1(out_cnt[4]), .I2(out_cnt[3]), .I3(out_cnt[2]), .O(n29897)
         );
  NR2 U25065 ( .I1(n29910), .I2(n30030), .O(n23599) );
  INV1S U25066 ( .I(n29967), .O(n23600) );
  OR2S U25067 ( .I1(n23600), .I2(n23770), .O(n23796) );
  INV1S U25068 ( .I(n23796), .O(n23814) );
  NR2 U25069 ( .I1(n23814), .I2(n16186), .O(n23832) );
  NR2 U25070 ( .I1(n23832), .I2(n30036), .O(n23620) );
  NR2 U25071 ( .I1(n23603), .I2(n23620), .O(n23821) );
  NR2 U25072 ( .I1(n23830), .I2(n23821), .O(n23829) );
  ND2S U25073 ( .I1(n23829), .I2(i_row[2]), .O(n23606) );
  XNR2HS U25074 ( .I1(i_row[2]), .I2(n23623), .O(n23602) );
  ND2S U25075 ( .I1(n23832), .I2(n23602), .O(n23605) );
  ND3S U25076 ( .I1(n23603), .I2(i_row[1]), .I3(n23827), .O(n23604) );
  ND3S U25077 ( .I1(n23606), .I2(n23605), .I3(n23604), .O(n13607) );
  NR3 U25078 ( .I1(n24025), .I2(n23607), .I3(n23730), .O(n23670) );
  NR2 U25079 ( .I1(n23675), .I2(n23670), .O(n23669) );
  ND2S U25080 ( .I1(n23669), .I2(n23900), .O(n23610) );
  ND2S U25081 ( .I1(n23675), .I2(img_size_hold[2]), .O(n23609) );
  INV1S U25082 ( .I(n23607), .O(n23611) );
  ND3S U25083 ( .I1(n30039), .I2(img_size[3]), .I3(n23611), .O(n23608) );
  ND3S U25084 ( .I1(n23610), .I2(n23609), .I3(n23608), .O(n13642) );
  ND2S U25085 ( .I1(n23669), .I2(img_size[3]), .O(n23614) );
  ND2S U25086 ( .I1(n23675), .I2(img_size_hold[3]), .O(n23613) );
  ND3S U25087 ( .I1(n30039), .I2(img_size[4]), .I3(n23611), .O(n23612) );
  ND3S U25088 ( .I1(n23614), .I2(n23613), .I3(n23612), .O(n13641) );
  AOI12HS U25089 ( .B1(n30018), .B2(n30014), .A1(addr[6]), .O(n23615) );
  AN2B1S U25090 ( .I1(n23616), .B1(n23615), .O(n13626) );
  NR2 U25091 ( .I1(rgb_value[23]), .I2(rgb_value[15]), .O(n29943) );
  INV1S U25092 ( .I(rgb_value[7]), .O(n29915) );
  ND2S U25093 ( .I1(n29943), .I2(n29915), .O(gray_max[7]) );
  ND2S U25094 ( .I1(n23682), .I2(n29910), .O(n31996) );
  ND2S U25095 ( .I1(n30030), .I2(n30032), .O(n29870) );
  NR3 U25096 ( .I1(out_cnt[2]), .I2(out_cnt[3]), .I3(n29870), .O(n23672) );
  ND2S U25097 ( .I1(n31997), .I2(n23672), .O(n23683) );
  XOR2HS U25098 ( .I1(n23683), .I2(out_cnt[4]), .O(n23617) );
  ND2S U25099 ( .I1(n23682), .I2(n23617), .O(n13682) );
  XOR3S U25100 ( .I1(rgb_value[14]), .I2(rgb_value[23]), .I3(rgb_value[7]), 
        .O(intadd_8_A_5_) );
  INV1S U25101 ( .I(temp_cnt[0]), .O(n29539) );
  AN4B1S U25102 ( .I1(n23619), .I2(n23618), .I3(n30007), .B1(addr[3]), .O(
        n23690) );
  NR2 U25103 ( .I1(n29539), .I2(n30019), .O(n23630) );
  ND2S U25104 ( .I1(temp_cnt[1]), .I2(n23630), .O(n23632) );
  ND2S U25105 ( .I1(n30021), .I2(n30019), .O(n23631) );
  OA112S U25106 ( .C1(temp_cnt[1]), .C2(n23630), .A1(n23632), .B1(n23631), .O(
        n13624) );
  ND2S U25107 ( .I1(n23620), .I2(n23622), .O(n23621) );
  MUX2S U25108 ( .A(n23622), .B(n23621), .S(i_row[1]), .O(n23627) );
  AN2S U25109 ( .I1(n23624), .I2(n23623), .O(n23625) );
  ND2S U25110 ( .I1(n23832), .I2(n23625), .O(n23626) );
  ND2S U25111 ( .I1(n23627), .I2(n23626), .O(n13608) );
  NR2 U25112 ( .I1(n29962), .I2(act_cnt[0]), .O(n23644) );
  ND2S U25113 ( .I1(n30036), .I2(n23640), .O(n23635) );
  NR2 U25114 ( .I1(n23644), .I2(n29961), .O(n29963) );
  ND2S U25115 ( .I1(n29964), .I2(in_valid2), .O(n29965) );
  AO12S U25116 ( .B1(n29963), .B2(n29965), .A1(n23649), .O(n23629) );
  ND2S U25117 ( .I1(n23629), .I2(n23628), .O(n13686) );
  INV1S U25118 ( .I(temp_cnt[2]), .O(n29542) );
  ND3S U25119 ( .I1(temp_cnt[1]), .I2(temp_cnt[2]), .I3(n23630), .O(n30024) );
  ND2S U25120 ( .I1(n30024), .I2(n23631), .O(n30022) );
  OAI22S U25121 ( .A1(n29542), .A2(n30022), .B1(n23632), .B2(n30022), .O(
        n13623) );
  INV1S U25122 ( .I(n29997), .O(n23633) );
  ND2S U25123 ( .I1(set_cnt[2]), .I2(n23633), .O(n30001) );
  AOI12HS U25124 ( .B1(set_cnt[2]), .B2(n29998), .A1(n23633), .O(n23634) );
  AN2B1S U25125 ( .I1(n30001), .B1(n23634), .O(n13635) );
  ND2S U25126 ( .I1(n23644), .I2(act_cnt[1]), .O(n23650) );
  OA12S U25127 ( .B1(n23650), .B2(act_cnt[2]), .A1(n23652), .O(n23656) );
  MUX2S U25128 ( .A(n23654), .B(act[16]), .S(n23656), .O(n13661) );
  ND2S U25129 ( .I1(n30039), .I2(act_ptr[0]), .O(n23638) );
  INV1S U25130 ( .I(n23638), .O(n23637) );
  ND2S U25131 ( .I1(n23638), .I2(n23635), .O(n23643) );
  INV1S U25132 ( .I(n23643), .O(n23636) );
  MUX2S U25133 ( .A(n23637), .B(n23636), .S(act_ptr[1]), .O(n13645) );
  OAI222S U25134 ( .A1(n23643), .A2(n23642), .B1(n23641), .B2(n23640), .C1(
        n23639), .C2(n23638), .O(n13684) );
  INV1S U25135 ( .I(n23644), .O(n23645) );
  NR2 U25136 ( .I1(act_cnt[1]), .I2(n23645), .O(n23647) );
  ND2S U25137 ( .I1(n23647), .I2(act_cnt[2]), .O(n23646) );
  ND2S U25138 ( .I1(n23646), .I2(n23652), .O(n23657) );
  MUX2S U25139 ( .A(act[10]), .B(n23654), .S(n23657), .O(n13667) );
  ND2S U25140 ( .I1(n23647), .I2(n23649), .O(n23648) );
  ND2S U25141 ( .I1(n23648), .I2(n23652), .O(n23660) );
  INV1S U25142 ( .I(act[22]), .O(n23885) );
  INV1S U25143 ( .I(n23648), .O(n23659) );
  MOAI1S U25144 ( .A1(n23660), .A2(n23885), .B1(n23659), .B2(action[1]), .O(
        n13655) );
  OA12S U25145 ( .B1(n23650), .B2(n23649), .A1(n23652), .O(n23658) );
  MUX2S U25146 ( .A(n23654), .B(act[4]), .S(n23658), .O(n13673) );
  ND2S U25147 ( .I1(n23651), .I2(act_cnt[2]), .O(n23653) );
  OA12S U25148 ( .B1(n23653), .B2(act_cnt[1]), .A1(n23652), .O(n23661) );
  MUX2S U25149 ( .A(n23654), .B(act[7]), .S(n23661), .O(n13670) );
  OA12S U25150 ( .B1(n23653), .B2(n29964), .A1(n23652), .O(n23662) );
  MUX2S U25151 ( .A(n23654), .B(act[1]), .S(n23662), .O(n13676) );
  MUX2S U25152 ( .A(n23655), .B(act[17]), .S(n23656), .O(n13662) );
  MUX2S U25153 ( .A(act[11]), .B(n23655), .S(n23657), .O(n13668) );
  INV1S U25154 ( .I(act[23]), .O(n23883) );
  MOAI1S U25155 ( .A1(n23660), .A2(n23883), .B1(n23659), .B2(action[2]), .O(
        n13656) );
  MUX2S U25156 ( .A(n23655), .B(act[5]), .S(n23658), .O(n13674) );
  MUX2S U25157 ( .A(n23655), .B(act[8]), .S(n23661), .O(n13671) );
  MUX2S U25158 ( .A(n23655), .B(act[2]), .S(n23662), .O(n13677) );
  MUX2S U25159 ( .A(n23663), .B(act[15]), .S(n23656), .O(n13663) );
  MUX2S U25160 ( .A(act[9]), .B(n23663), .S(n23657), .O(n13669) );
  MUX2S U25161 ( .A(n23663), .B(act[3]), .S(n23658), .O(n13675) );
  MOAI1S U25162 ( .A1(n23660), .A2(n23884), .B1(n23659), .B2(action[0]), .O(
        n13657) );
  MUX2S U25163 ( .A(n23663), .B(act[6]), .S(n23661), .O(n13672) );
  MUX2S U25164 ( .A(n23663), .B(act[0]), .S(n23662), .O(n13678) );
  OR2S U25165 ( .I1(image_size[0]), .I2(n23666), .O(n23668) );
  MOAI1S U25166 ( .A1(n23668), .A2(image_size[1]), .B1(img_size_hold[2]), .B2(
        n23666), .O(n11201) );
  INV1S U25167 ( .I(image_size[1]), .O(n23667) );
  MOAI1S U25168 ( .A1(n23667), .A2(n23664), .B1(n23666), .B2(img_size_hold[5]), 
        .O(n11204) );
  INV1S U25169 ( .I(n23669), .O(n23671) );
  MOAI1S U25170 ( .A1(n23671), .A2(n23665), .B1(n23675), .B2(img_size_hold[5]), 
        .O(n13639) );
  MOAI1S U25171 ( .A1(n23668), .A2(n23667), .B1(img_size_hold[4]), .B2(n23666), 
        .O(n11203) );
  AO222S U25172 ( .A1(img_size[4]), .A2(n23669), .B1(n23670), .B2(img_size[5]), 
        .C1(n23675), .C2(img_size_hold[4]), .O(n13640) );
  INV1S U25173 ( .I(img_size[1]), .O(n24030) );
  MOAI1S U25174 ( .A1(n23671), .A2(n24030), .B1(n23900), .B2(n23670), .O(
        n13643) );
  MOAI1S U25175 ( .A1(n23671), .A2(n28540), .B1(img_size[1]), .B2(n23670), .O(
        n13689) );
  INV1S U25176 ( .I(out_cnt[2]), .O(n29793) );
  MOAI1S U25177 ( .A1(n29793), .A2(n29870), .B1(n29793), .B2(n29870), .O(
        n23676) );
  ND2S U25178 ( .I1(n23672), .I2(n30033), .O(n23673) );
  ND2S U25179 ( .I1(n31997), .I2(n23673), .O(n23677) );
  ND2S U25180 ( .I1(n29910), .I2(out_cnt[2]), .O(n23674) );
  OAI22S U25181 ( .A1(n23676), .A2(n23677), .B1(n23675), .B2(n23674), .O(
        n13680) );
  NR2 U25182 ( .I1(out_cnt[2]), .I2(n29870), .O(n23678) );
  MOAI1S U25183 ( .A1(n23678), .A2(n23677), .B1(n29910), .B2(n23682), .O(
        n23679) );
  MOAI1S U25184 ( .A1(n23683), .A2(n30033), .B1(n23679), .B2(out_cnt[3]), .O(
        n13679) );
  NR2 U25185 ( .I1(out_cnt[0]), .I2(n29910), .O(n23680) );
  XNR2HS U25186 ( .I1(n23680), .I2(out_cnt[1]), .O(n23681) );
  OAI112HS U25187 ( .C1(out_cnt[4]), .C2(n23683), .A1(n23682), .B1(n23681), 
        .O(n13683) );
  INV1S U25188 ( .I(col[3]), .O(n24228) );
  INV1S U25189 ( .I(col[2]), .O(n23905) );
  INV1S U25190 ( .I(col[1]), .O(n23732) );
  ND2S U25191 ( .I1(n23740), .I2(col[1]), .O(n23685) );
  NR2 U25192 ( .I1(n28555), .I2(col[0]), .O(n23684) );
  AOI22S U25193 ( .A1(n23870), .A2(n23732), .B1(n23685), .B2(n23684), .O(
        n23687) );
  ND2S U25194 ( .I1(n23791), .I2(n23905), .O(n23686) );
  MOAI1S U25195 ( .A1(n23791), .A2(n23905), .B1(n23687), .B2(n23686), .O(
        n23689) );
  ND2S U25196 ( .I1(n23795), .I2(n24228), .O(n23688) );
  MOAI1S U25197 ( .A1(n23795), .A2(n24228), .B1(n23689), .B2(n23688), .O(
        n23697) );
  INV1S U25198 ( .I(n23797), .O(n23696) );
  OAI12HS U25199 ( .B1(c_s[0]), .B2(n23694), .A1(n23693), .O(n24705) );
  INV1S U25200 ( .I(n24705), .O(n23695) );
  ND3S U25201 ( .I1(n23697), .I2(n23696), .I3(n23695), .O(n23710) );
  OA12S U25202 ( .B1(n23698), .B2(img_size[4]), .A1(img_size[5]), .O(n23700)
         );
  NR2 U25203 ( .I1(n23700), .I2(n23699), .O(n23766) );
  INV1S U25204 ( .I(n23701), .O(n23702) );
  NR2 U25205 ( .I1(n23702), .I2(n24031), .O(n23747) );
  OR2S U25206 ( .I1(col[1]), .I2(n23747), .O(n23705) );
  NR2 U25207 ( .I1(col[2]), .I2(n23749), .O(n23704) );
  NR2 U25208 ( .I1(col[3]), .I2(n23751), .O(n23703) );
  NR2 U25209 ( .I1(n23704), .I2(n23703), .O(n23707) );
  OAI112HS U25210 ( .C1(img_size[1]), .C2(col[0]), .A1(n23705), .B1(n23707), 
        .O(n23759) );
  INV1S U25211 ( .I(n23749), .O(n23706) );
  MOAI1S U25212 ( .A1(n23905), .A2(n23706), .B1(col[1]), .B2(n23747), .O(
        n23760) );
  ND2S U25213 ( .I1(n23707), .I2(n23760), .O(n23708) );
  ND2S U25214 ( .I1(n23751), .I2(col[3]), .O(n23762) );
  ND3S U25215 ( .I1(n23759), .I2(n23708), .I3(n23762), .O(n23709) );
  MOAI1S U25216 ( .A1(n23812), .A2(n23710), .B1(n23766), .B2(n23709), .O(
        n23721) );
  XNR2HS U25217 ( .I1(img_size[3]), .I2(n23954), .O(n23867) );
  INV1S U25218 ( .I(cal_cnt[4]), .O(n23716) );
  AOI22S U25219 ( .A1(cal_cnt[3]), .A2(n23869), .B1(n23867), .B2(cal_cnt[4]), 
        .O(n23715) );
  INV1S U25220 ( .I(cal_cnt[2]), .O(n29973) );
  NR2 U25221 ( .I1(cal_cnt[2]), .I2(n24030), .O(n23712) );
  ND2S U25222 ( .I1(n28555), .I2(cal_cnt[1]), .O(n23711) );
  OAI22S U25223 ( .A1(n29973), .A2(n23870), .B1(n23712), .B2(n23711), .O(
        n23713) );
  OAI12HS U25224 ( .B1(cal_cnt[3]), .B2(n23869), .A1(n23713), .O(n23714) );
  AOI22S U25225 ( .A1(n23795), .A2(n23716), .B1(n23715), .B2(n23714), .O(
        n23720) );
  NR3 U25226 ( .I1(cal_cnt[5]), .I2(cal_cnt[6]), .I3(cal_cnt[8]), .O(n23718)
         );
  INV1S U25227 ( .I(cal_cnt[7]), .O(n23717) );
  OAI12HS U25228 ( .B1(n23720), .B2(n23719), .A1(n23770), .O(n23901) );
  AN3B2S U25229 ( .I1(n23901), .B1(n23812), .B2(n24705), .O(n23737) );
  NR2 U25230 ( .I1(n23721), .I2(n23737), .O(n23729) );
  XNR2HS U25231 ( .I1(col[3]), .I2(n23867), .O(n23722) );
  NR2 U25232 ( .I1(n23722), .I2(n23797), .O(n23728) );
  XNR2HS U25233 ( .I1(col[2]), .I2(n23869), .O(n23726) );
  XOR2HS U25234 ( .I1(col[1]), .I2(n23740), .O(n23724) );
  XOR2HS U25235 ( .I1(col[0]), .I2(n28555), .O(n23723) );
  ND2S U25236 ( .I1(n23724), .I2(n23723), .O(n23725) );
  NR2 U25237 ( .I1(n23726), .I2(n23725), .O(n23727) );
  AN2S U25238 ( .I1(n23728), .I2(n23727), .O(n23771) );
  ND2S U25239 ( .I1(n23771), .I2(n24705), .O(n23774) );
  INV1S U25240 ( .I(n23739), .O(n23731) );
  MUX2S U25241 ( .A(n23731), .B(n23737), .S(col[0]), .O(n13615) );
  NR2 U25242 ( .I1(col[0]), .I2(n23732), .O(n24015) );
  INV1S U25243 ( .I(col[0]), .O(n23763) );
  NR2 U25244 ( .I1(col[1]), .I2(n23763), .O(n24019) );
  NR2 U25245 ( .I1(n24015), .I2(n24019), .O(n23733) );
  MOAI1S U25246 ( .A1(n23739), .A2(n23733), .B1(col[1]), .B2(n23737), .O(
        n13621) );
  INV1S U25247 ( .I(n23737), .O(n23736) );
  NR2 U25248 ( .I1(n23905), .I2(n24147), .O(n24226) );
  NR2 U25249 ( .I1(n24226), .I2(n23739), .O(n23735) );
  ND2S U25250 ( .I1(n24147), .I2(n23905), .O(n23734) );
  MOAI1S U25251 ( .A1(n23736), .A2(n23905), .B1(n23735), .B2(n23734), .O(
        n13614) );
  XOR2HS U25252 ( .I1(n24228), .I2(n24226), .O(n23738) );
  MOAI1S U25253 ( .A1(n23739), .A2(n23738), .B1(col[3]), .B2(n23737), .O(
        n13620) );
  XNR2HS U25254 ( .I1(row[2]), .I2(n23869), .O(n23744) );
  XOR2HS U25255 ( .I1(row[1]), .I2(n23740), .O(n23742) );
  XOR2HS U25256 ( .I1(row[0]), .I2(n28555), .O(n23741) );
  ND2S U25257 ( .I1(n23742), .I2(n23741), .O(n23743) );
  NR2 U25258 ( .I1(n23744), .I2(n23743), .O(n23745) );
  ND2S U25259 ( .I1(n13942), .I2(n23745), .O(n23769) );
  INV1S U25260 ( .I(row[0]), .O(n23776) );
  ND2S U25261 ( .I1(n23776), .I2(n24030), .O(n23746) );
  FA1S U25262 ( .A(row[1]), .B(n23747), .CI(n23746), .CO(n23748) );
  FA1S U25263 ( .A(n23749), .B(row[2]), .CI(n23748), .CO(n23750) );
  MAO222S U25264 ( .A1(row[3]), .B1(n23751), .C1(n23750), .O(n23767) );
  INV1S U25265 ( .I(row[1]), .O(n23775) );
  NR2 U25266 ( .I1(n23775), .I2(n23870), .O(n23753) );
  OR2S U25267 ( .I1(n28555), .I2(row[0]), .O(n23752) );
  MOAI1S U25268 ( .A1(n23753), .A2(n23752), .B1(n23870), .B2(n23775), .O(
        n23755) );
  NR2 U25269 ( .I1(row[2]), .I2(n23869), .O(n23754) );
  INV1S U25270 ( .I(row[2]), .O(n24010) );
  OAI22S U25271 ( .A1(n23755), .A2(n23754), .B1(n23791), .B2(n24010), .O(
        n23757) );
  INV1S U25272 ( .I(row[3]), .O(n24011) );
  ND2S U25273 ( .I1(n23795), .I2(n24011), .O(n23756) );
  INV1S U25274 ( .I(n23759), .O(n23765) );
  INV1S U25275 ( .I(n23760), .O(n23761) );
  ND3S U25276 ( .I1(n23766), .I2(n23765), .I3(n23764), .O(n23772) );
  MXL2HS U25277 ( .A(n23767), .B(n23758), .S(n23772), .OB(n23768) );
  MXL2HS U25278 ( .A(n23769), .B(n23768), .S(n23774), .OB(n23781) );
  ND2S U25279 ( .I1(n23771), .I2(n23770), .O(n23773) );
  INV1S U25280 ( .I(n23783), .O(n23777) );
  NR2 U25281 ( .I1(n23781), .I2(n23777), .O(n23780) );
  MUX2S U25282 ( .A(n23780), .B(n23777), .S(row[0]), .O(n13619) );
  INV1S U25283 ( .I(n23780), .O(n23779) );
  NR2 U25284 ( .I1(row[0]), .I2(n23775), .O(n23914) );
  NR2 U25285 ( .I1(row[1]), .I2(n23776), .O(n23967) );
  NR2 U25286 ( .I1(n23914), .I2(n23967), .O(n23778) );
  MOAI1S U25287 ( .A1(n23779), .A2(n23778), .B1(row[1]), .B2(n23777), .O(
        n13616) );
  INV1S U25288 ( .I(n24099), .O(n23908) );
  ND2S U25289 ( .I1(n23780), .I2(n23908), .O(n23787) );
  INV1S U25290 ( .I(n23787), .O(n23785) );
  INV1S U25291 ( .I(n23781), .O(n23782) );
  OAI12HS U25292 ( .B1(n24010), .B2(n24099), .A1(n23782), .O(n23784) );
  ND2S U25293 ( .I1(n23784), .I2(n23783), .O(n23786) );
  OA12S U25294 ( .B1(n23785), .B2(row[2]), .A1(n23786), .O(n13617) );
  MOAI1S U25295 ( .A1(n23787), .A2(n24098), .B1(row[3]), .B2(n23786), .O(
        n13618) );
  NR2 U25296 ( .I1(n28555), .I2(i_col[0]), .O(n23789) );
  FA1S U25297 ( .A(n23870), .B(n23789), .CI(n23788), .CO(n23790) );
  FA1S U25298 ( .A(n23792), .B(n23791), .CI(n23790), .CO(n23793) );
  MAO222S U25299 ( .A1(n23795), .B1(n23794), .C1(n23793), .O(n23798) );
  OAI12HS U25300 ( .B1(n23798), .B2(n23797), .A1(n23796), .O(n23799) );
  NR2 U25301 ( .I1(n23799), .I2(n30039), .O(n23820) );
  ND2S U25302 ( .I1(n23801), .I2(n23800), .O(n23802) );
  ND2S U25303 ( .I1(n23803), .I2(n23802), .O(n23806) );
  AOI13HS U25304 ( .B1(n23807), .B2(n23806), .B3(n23805), .A1(n23804), .O(
        n23809) );
  ND2P U25305 ( .I1(n23808), .I2(n23812), .O(n23850) );
  NR2 U25306 ( .I1(n23809), .I2(n23850), .O(n23810) );
  AO12S U25307 ( .B1(i_col[0]), .B2(n23820), .A1(n23810), .O(n23833) );
  ND2S U25308 ( .I1(n23833), .I2(i_col[1]), .O(n23837) );
  INV1S U25309 ( .I(n23837), .O(n23816) );
  INV1S U25310 ( .I(n23810), .O(n23818) );
  ND2S U25311 ( .I1(n23811), .I2(n23820), .O(n23815) );
  INV1S U25312 ( .I(n23812), .O(n23813) );
  ND2S U25313 ( .I1(n23814), .I2(n23813), .O(n23817) );
  OAI112HS U25314 ( .C1(i_col[1]), .C2(n23818), .A1(n23815), .B1(n23817), .O(
        n23836) );
  MUX2S U25315 ( .A(n23816), .B(n23836), .S(i_col[2]), .O(n13611) );
  ND2S U25316 ( .I1(n23818), .I2(n23817), .O(n23819) );
  MUX2S U25317 ( .A(n23820), .B(n23819), .S(i_col[0]), .O(n13613) );
  INV1S U25318 ( .I(n23821), .O(n23822) );
  MUX2S U25319 ( .A(n23832), .B(n23822), .S(i_row[0]), .O(n13609) );
  ND2S U25320 ( .I1(n23823), .I2(i_row[0]), .O(n23826) );
  OAI12HS U25321 ( .B1(n23827), .B2(n23824), .A1(n23828), .O(n23825) );
  MUX2S U25322 ( .A(n23830), .B(n23829), .S(n23828), .O(n23831) );
  AO12S U25323 ( .B1(n23832), .B2(n13941), .A1(n23831), .O(n13606) );
  OA12S U25324 ( .B1(i_col[1]), .B2(n23833), .A1(n23836), .O(n13610) );
  NR2 U25325 ( .I1(n23835), .I2(n23834), .O(n23838) );
  MOAI1S U25326 ( .A1(n23838), .A2(n23837), .B1(n23836), .B2(i_col[3]), .O(
        n13612) );
  INV1S U25327 ( .I(n23840), .O(n23842) );
  NR2P U25328 ( .I1(n23842), .I2(n23841), .O(n28534) );
  ND2 U25329 ( .I1(n23844), .I2(n23843), .O(n28529) );
  OAI22S U25330 ( .A1(n23846), .A2(n28530), .B1(n13897), .B2(n23845), .O(
        n23847) );
  OAI12HS U25331 ( .B1(n28536), .B2(n21504), .A1(n23849), .O(n23892) );
  NR2F U25332 ( .I1(n24025), .I2(n23850), .O(n28575) );
  INV1S U25333 ( .I(n23851), .O(n23854) );
  INV1S U25334 ( .I(n29968), .O(n23853) );
  INV1S U25335 ( .I(n23894), .O(n24706) );
  INV1S U25336 ( .I(n23900), .O(n23855) );
  NR2 U25337 ( .I1(n23856), .I2(n23870), .O(n28552) );
  NR2 U25338 ( .I1(n23857), .I2(n23870), .O(n28551) );
  NR2 U25339 ( .I1(n23858), .I2(n23870), .O(n28550) );
  ND2S U25340 ( .I1(n28550), .I2(A67_shift[79]), .O(n23864) );
  INV1S U25341 ( .I(n23859), .O(n23861) );
  NR2 U25342 ( .I1(n28540), .I2(n23860), .O(n23929) );
  NR2 U25343 ( .I1(n23929), .I2(n23954), .O(n23868) );
  NR2 U25344 ( .I1(n23861), .I2(n23868), .O(n28554) );
  NR2 U25345 ( .I1(n23862), .I2(n23870), .O(n28553) );
  AOI22S U25346 ( .A1(A67_shift[111]), .A2(n28554), .B1(A67_shift[15]), .B2(
        n28553), .O(n23863) );
  NR2 U25347 ( .I1(n23866), .I2(n23865), .O(n23873) );
  NR2 U25348 ( .I1(n23868), .I2(n23867), .O(n28547) );
  INV1S U25349 ( .I(n26653), .O(n28546) );
  INV1S U25350 ( .I(n28544), .O(n28545) );
  AOI22S U25351 ( .A1(n28546), .A2(A67_shift[175]), .B1(n28545), .B2(
        A67_shift[47]), .O(n23871) );
  ND2S U25352 ( .I1(n28550), .I2(A67_shift[95]), .O(n23875) );
  AOI22S U25353 ( .A1(n28554), .A2(A67_shift[127]), .B1(n28551), .B2(
        A67_shift[223]), .O(n23874) );
  NR2 U25354 ( .I1(n23877), .I2(n23876), .O(n23880) );
  AOI22S U25355 ( .A1(n28546), .A2(A67_shift[191]), .B1(n28545), .B2(
        A67_shift[63]), .O(n23878) );
  NR2 U25356 ( .I1(act[22]), .I2(n23884), .O(n28564) );
  ND2S U25357 ( .I1(n28564), .I2(gray_avg_out[7]), .O(n23888) );
  NR2 U25358 ( .I1(act[21]), .I2(n23885), .O(n28565) );
  ND2S U25359 ( .I1(n28565), .I2(gray_weight_out[7]), .O(n23887) );
  NR2 U25360 ( .I1(act[21]), .I2(act[22]), .O(n28566) );
  ND2S U25361 ( .I1(n28566), .I2(gray_max_out[7]), .O(n23886) );
  AOI12HT U25362 ( .B1(n23892), .B2(n28575), .A1(n23891), .O(n24581) );
  INV1S U25363 ( .I(n23895), .O(n23893) );
  AOI22S U25364 ( .A1(n13773), .A2(img[591]), .B1(n29407), .B2(n30037), .O(
        n23896) );
  ND2S U25365 ( .I1(n24340), .I2(n23896), .O(n23903) );
  NR2 U25366 ( .I1(col[2]), .I2(n24228), .O(n24014) );
  INV1S U25367 ( .I(n24014), .O(n24220) );
  INV1S U25368 ( .I(n24019), .O(n24022) );
  NR2 U25369 ( .I1(n24220), .I2(n24022), .O(n23899) );
  NR2 U25370 ( .I1(n23899), .I2(n24692), .O(n24105) );
  NR2 U25371 ( .I1(n23901), .I2(n30039), .O(n24702) );
  OR2T U25372 ( .I1(n24702), .I2(n13908), .O(n24012) );
  NR2 U25373 ( .I1(n24002), .I2(n24099), .O(n24640) );
  OR2 U25374 ( .I1(n24640), .I2(n24692), .O(n24689) );
  NR2P U25375 ( .I1(n24240), .I2(n24689), .O(n24693) );
  AO12 U25376 ( .B1(n24105), .B2(n24694), .A1(n24693), .O(n28578) );
  MUX2 U25377 ( .A(n23903), .B(img[567]), .S(n28578), .O(n12971) );
  AOI22S U25378 ( .A1(n13773), .A2(img[567]), .B1(n13779), .B2(n30038), .O(
        n23904) );
  ND2S U25379 ( .I1(n24340), .I2(n23904), .O(n23906) );
  NR2 U25380 ( .I1(col[3]), .I2(n23905), .O(n24152) );
  NR2 U25381 ( .I1(n24134), .I2(n24692), .O(n24006) );
  AO12 U25382 ( .B1(n24006), .B2(n24694), .A1(n24693), .O(n28581) );
  MUX2 U25383 ( .A(n23906), .B(img[591]), .S(n28581), .O(n12941) );
  AOI22S U25384 ( .A1(n13773), .A2(img[79]), .B1(n29242), .B2(n30040), .O(
        n23907) );
  ND2S U25385 ( .I1(n24340), .I2(n23907), .O(n23910) );
  NR2 U25386 ( .I1(n24011), .I2(n24010), .O(n23974) );
  MUX2 U25387 ( .A(img[55]), .B(n23910), .S(n28584), .O(n13480) );
  AOI22S U25388 ( .A1(n13773), .A2(img[55]), .B1(n27049), .B2(n30041), .O(
        n23911) );
  ND2S U25389 ( .I1(n24340), .I2(n23911), .O(n23912) );
  AOI22S U25390 ( .A1(n13780), .A2(img[1271]), .B1(n29407), .B2(n30042), .O(
        n23913) );
  ND2S U25391 ( .I1(n24340), .I2(n23913), .O(n23917) );
  INV1S U25392 ( .I(n23914), .O(n24051) );
  INV1S U25393 ( .I(n23961), .O(n23915) );
  NR2 U25394 ( .I1(n28540), .I2(n24495), .O(n24614) );
  NR2 U25395 ( .I1(n24463), .I2(n24726), .O(n23916) );
  INV1S U25396 ( .I(n24015), .O(n24029) );
  NR2 U25397 ( .I1(n24139), .I2(n24029), .O(n24766) );
  MUX2 U25398 ( .A(img[1167]), .B(n23917), .S(n28590), .O(n12371) );
  AOI22S U25399 ( .A1(n28862), .A2(n30043), .B1(n27919), .B2(img[1167]), .O(
        n23921) );
  ND3S U25400 ( .I1(n24340), .I2(n23921), .I3(n23920), .O(n23930) );
  NR2 U25401 ( .I1(n24234), .I2(n24022), .O(n24670) );
  NR2 U25402 ( .I1(img_size[3]), .I2(n24698), .O(n23924) );
  INV1S U25403 ( .I(n23924), .O(n23928) );
  NR2 U25404 ( .I1(n23922), .I2(n23928), .O(n23927) );
  INV1S U25405 ( .I(n23923), .O(n23925) );
  OAI12HS U25406 ( .B1(n24700), .B2(n23925), .A1(n24033), .O(n24541) );
  MUX2 U25407 ( .A(img[1271]), .B(n23930), .S(n28595), .O(n12261) );
  AOI22S U25408 ( .A1(n26970), .A2(img[1231]), .B1(n29397), .B2(n30044), .O(
        n23931) );
  ND2S U25409 ( .I1(n24340), .I2(n23931), .O(n23934) );
  NR2P U25410 ( .I1(n24463), .I2(n24692), .O(n24466) );
  NR3 U25411 ( .I1(n23932), .I2(n24030), .I3(n24699), .O(n23933) );
  NR2P U25412 ( .I1(n23933), .I2(n24240), .O(n24748) );
  AOI22S U25413 ( .A1(n29242), .A2(n30045), .B1(n27919), .B2(img[1207]), .O(
        n23936) );
  ND2S U25414 ( .I1(n13770), .I2(img[1271]), .O(n23935) );
  ND3S U25415 ( .I1(n24340), .I2(n23936), .I3(n23935), .O(n23937) );
  MUX2 U25416 ( .A(img[1231]), .B(n23937), .S(n28602), .O(n12307) );
  AOI22S U25417 ( .A1(n13778), .A2(img[1399]), .B1(n25859), .B2(n30046), .O(
        n23938) );
  ND2S U25418 ( .I1(n24340), .I2(n23938), .O(n23940) );
  INV1S U25419 ( .I(n23967), .O(n24013) );
  NR2 U25420 ( .I1(n24726), .I2(n24476), .O(n23939) );
  AOI22S U25421 ( .A1(n25591), .A2(n30047), .B1(n24313), .B2(img[1295]), .O(
        n23943) );
  ND2S U25422 ( .I1(n13902), .I2(img[1359]), .O(n23942) );
  ND3S U25423 ( .I1(n24340), .I2(n23943), .I3(n23942), .O(n23944) );
  MUX2 U25424 ( .A(img[1399]), .B(n23944), .S(n28609), .O(n12139) );
  AOI22S U25425 ( .A1(n26822), .A2(img[1359]), .B1(n29397), .B2(n30048), .O(
        n23945) );
  ND2S U25426 ( .I1(n24340), .I2(n23945), .O(n23946) );
  MUX2 U25427 ( .A(n23946), .B(img[1335]), .S(n28612), .O(n12203) );
  AOI22S U25428 ( .A1(n27735), .A2(n30049), .B1(n27919), .B2(img[1335]), .O(
        n23948) );
  ND3S U25429 ( .I1(n24340), .I2(n23948), .I3(n23947), .O(n23949) );
  MUX2 U25430 ( .A(img[1359]), .B(n23949), .S(n28617), .O(n12173) );
  AOI22S U25431 ( .A1(n27065), .A2(img[975]), .B1(n28862), .B2(n30050), .O(
        n23950) );
  ND2S U25432 ( .I1(n24340), .I2(n23950), .O(n23952) );
  NR2 U25433 ( .I1(n24002), .I2(n24112), .O(n24646) );
  ND2S U25434 ( .I1(n24748), .I2(n24713), .O(n23951) );
  AOI22S U25435 ( .A1(n28106), .A2(img[951]), .B1(n28862), .B2(n30051), .O(
        n23953) );
  ND2S U25436 ( .I1(n24340), .I2(n23953), .O(n23959) );
  INV1S U25437 ( .I(n23954), .O(n23955) );
  NR2 U25438 ( .I1(n24698), .I2(n23955), .O(n23957) );
  OAI12HS U25439 ( .B1(n24033), .B2(n23957), .A1(n23956), .O(n24716) );
  NR2 U25440 ( .I1(n24134), .I2(n24716), .O(n23958) );
  NR2P U25441 ( .I1(n24646), .I2(n24716), .O(n24717) );
  NR2P U25442 ( .I1(n23958), .I2(n24717), .O(n28623) );
  MUX2 U25443 ( .A(img[975]), .B(n23959), .S(n28623), .O(n12563) );
  AOI22S U25444 ( .A1(n28347), .A2(img[207]), .B1(n27511), .B2(n30052), .O(
        n23960) );
  ND2S U25445 ( .I1(n24340), .I2(n23960), .O(n23963) );
  INV1S U25446 ( .I(n24105), .O(n23962) );
  MUX2 U25447 ( .A(img[183]), .B(n23963), .S(n28626), .O(n13349) );
  AOI22S U25448 ( .A1(n26970), .A2(img[183]), .B1(n13775), .B2(n30053), .O(
        n23964) );
  ND2S U25449 ( .I1(n24340), .I2(n23964), .O(n23965) );
  MUX2 U25450 ( .A(img[207]), .B(n23965), .S(n28629), .O(n13331) );
  AOI22S U25451 ( .A1(n27957), .A2(img[335]), .B1(n28037), .B2(n30054), .O(
        n23966) );
  ND2S U25452 ( .I1(n24340), .I2(n23966), .O(n23969) );
  OAI12HS U25453 ( .B1(n24732), .B2(n24105), .A1(n24495), .O(n28632) );
  MUX2 U25454 ( .A(img[311]), .B(n23969), .S(n28632), .O(n13227) );
  AOI22S U25455 ( .A1(n13776), .A2(img[311]), .B1(n13775), .B2(n30055), .O(
        n23970) );
  ND2S U25456 ( .I1(n24340), .I2(n23970), .O(n23971) );
  OAI12HS U25457 ( .B1(n24732), .B2(n24006), .A1(n24495), .O(n28635) );
  AOI22S U25458 ( .A1(n26970), .A2(img[463]), .B1(n23918), .B2(n30056), .O(
        n23972) );
  ND2S U25459 ( .I1(n24340), .I2(n23972), .O(n23977) );
  ND2 U25460 ( .I1(n24203), .I2(n24664), .O(n24668) );
  INV1S U25461 ( .I(n23975), .O(n24741) );
  ND2S U25462 ( .I1(n24741), .I2(n24105), .O(n23976) );
  ND2S U25463 ( .I1(n24668), .I2(n23976), .O(n28638) );
  MUX2 U25464 ( .A(n23977), .B(img[439]), .S(n28638), .O(n13093) );
  AOI22S U25465 ( .A1(n13773), .A2(img[439]), .B1(n28182), .B2(n30057), .O(
        n23978) );
  ND2S U25466 ( .I1(n24340), .I2(n23978), .O(n23980) );
  ND2S U25467 ( .I1(n24741), .I2(n24006), .O(n23979) );
  ND2S U25468 ( .I1(n24668), .I2(n23979), .O(n28641) );
  AOI22S U25469 ( .A1(n13773), .A2(img[1527]), .B1(n28343), .B2(n30058), .O(
        n23981) );
  ND2S U25470 ( .I1(n24340), .I2(n23981), .O(n23984) );
  INV1S U25471 ( .I(n23982), .O(n23983) );
  INV1S U25472 ( .I(n24515), .O(n24509) );
  MUX2 U25473 ( .A(n23984), .B(img[1423]), .S(n28645), .O(n12115) );
  AOI22S U25474 ( .A1(n25377), .A2(n30059), .B1(n24946), .B2(img[1423]), .O(
        n23986) );
  ND3S U25475 ( .I1(n24340), .I2(n23986), .I3(n23985), .O(n23988) );
  AOI22S U25476 ( .A1(n13773), .A2(img[1487]), .B1(n28135), .B2(n30060), .O(
        n23989) );
  ND2S U25477 ( .I1(n24340), .I2(n23989), .O(n23990) );
  AOI22S U25478 ( .A1(n28162), .A2(n30061), .B1(n25444), .B2(img[1463]), .O(
        n23992) );
  ND2S U25479 ( .I1(n29124), .I2(img[1527]), .O(n23991) );
  ND3S U25480 ( .I1(n24340), .I2(n23992), .I3(n23991), .O(n23993) );
  MUX2 U25481 ( .A(img[1487]), .B(n23993), .S(n28656), .O(n12051) );
  AOI22S U25482 ( .A1(n13773), .A2(img[847]), .B1(n25859), .B2(n30062), .O(
        n23994) );
  ND2S U25483 ( .I1(n24340), .I2(n23994), .O(n23995) );
  INV1S U25484 ( .I(img[847]), .O(n23996) );
  AOI22S U25485 ( .A1(n13773), .A2(img[823]), .B1(n25377), .B2(n23996), .O(
        n23997) );
  ND2S U25486 ( .I1(n24340), .I2(n23997), .O(n23999) );
  ND2S U25487 ( .I1(n24748), .I2(n24006), .O(n23998) );
  AOI22S U25488 ( .A1(n13773), .A2(img[719]), .B1(n28862), .B2(n30063), .O(
        n24000) );
  ND2S U25489 ( .I1(n24340), .I2(n24000), .O(n24004) );
  NR2 U25490 ( .I1(n26653), .I2(n24699), .O(n24001) );
  NR2P U25491 ( .I1(n24001), .I2(n24240), .O(n24758) );
  NR2 U25492 ( .I1(n24002), .I2(n24051), .O(n24681) );
  ND2P U25493 ( .I1(n24758), .I2(n24753), .O(n24760) );
  ND2S U25494 ( .I1(n24758), .I2(n24105), .O(n24003) );
  AOI22S U25495 ( .A1(n13773), .A2(img[695]), .B1(n28162), .B2(n30064), .O(
        n24005) );
  ND2S U25496 ( .I1(n24340), .I2(n24005), .O(n24008) );
  ND2S U25497 ( .I1(n24758), .I2(n24006), .O(n24007) );
  AOI22S U25498 ( .A1(n13778), .A2(img[1879]), .B1(n13781), .B2(n30065), .O(
        n24009) );
  ND2S U25499 ( .I1(n24340), .I2(n24009), .O(n24016) );
  ND3P U25500 ( .I1(n24012), .I2(n24011), .I3(n24010), .O(n24111) );
  NR2 U25501 ( .I1(n24568), .I2(n24692), .O(n24563) );
  MUX2 U25502 ( .A(n24016), .B(img[1839]), .S(n28672), .O(n11693) );
  AOI22S U25503 ( .A1(n25377), .A2(n30066), .B1(n25444), .B2(img[1839]), .O(
        n24018) );
  ND3S U25504 ( .I1(n24340), .I2(n24018), .I3(n24017), .O(n24020) );
  MUX2 U25505 ( .A(img[1879]), .B(n24020), .S(n28676), .O(n11659) );
  AOI22S U25506 ( .A1(n26822), .A2(img[1903]), .B1(n28938), .B2(n30067), .O(
        n24021) );
  ND2S U25507 ( .I1(n24340), .I2(n24021), .O(n24024) );
  NR2 U25508 ( .I1(n24139), .I2(n24022), .O(n24490) );
  NR2 U25509 ( .I1(n24490), .I2(n24692), .O(n24023) );
  MUX2 U25510 ( .A(n24024), .B(img[1815]), .S(n28679), .O(n11723) );
  AOI22S U25511 ( .A1(n28938), .A2(n30068), .B1(n25444), .B2(img[1815]), .O(
        n24028) );
  INV1S U25512 ( .I(n24025), .O(n24026) );
  NR2 U25513 ( .I1(n24026), .I2(n24700), .O(n28908) );
  AOI22S U25514 ( .A1(n13903), .A2(img[1879]), .B1(img[1911]), .B2(n13782), 
        .O(n24027) );
  ND3S U25515 ( .I1(n24340), .I2(n24028), .I3(n24027), .O(n24036) );
  NR2 U25516 ( .I1(n24234), .I2(n24029), .O(n24542) );
  NR2 U25517 ( .I1(n28540), .I2(n24030), .O(n24035) );
  INV1S U25518 ( .I(n24031), .O(n24032) );
  MUX2 U25519 ( .A(img[1903]), .B(n24036), .S(n28683), .O(n11629) );
  AOI22S U25520 ( .A1(n29435), .A2(img[1911]), .B1(n13775), .B2(n30069), .O(
        n24037) );
  ND2S U25521 ( .I1(n24340), .I2(n24037), .O(n24039) );
  NR2 U25522 ( .I1(n24726), .I2(n24250), .O(n24038) );
  BUF12CK U25523 ( .I(n24581), .O(n24340) );
  AOI22S U25524 ( .A1(n28938), .A2(n30070), .B1(n27919), .B2(img[1807]), .O(
        n24041) );
  AOI22S U25525 ( .A1(n13905), .A2(img[1871]), .B1(img[1903]), .B2(n13782), 
        .O(n24040) );
  ND3S U25526 ( .I1(n24340), .I2(n24041), .I3(n24040), .O(n24044) );
  OAI12HS U25527 ( .B1(n24699), .B2(n24043), .A1(n24042), .O(n24235) );
  MUX2 U25528 ( .A(img[1911]), .B(n24044), .S(n28690), .O(n11627) );
  AOI22S U25529 ( .A1(n28318), .A2(img[1871]), .B1(n24374), .B2(n30071), .O(
        n24045) );
  ND2S U25530 ( .I1(n24340), .I2(n24045), .O(n24046) );
  AOI22S U25531 ( .A1(n28913), .A2(n30072), .B1(n24313), .B2(img[1847]), .O(
        n24048) );
  ND2S U25532 ( .I1(n13903), .I2(img[1911]), .O(n24047) );
  ND3S U25533 ( .I1(n24340), .I2(n24048), .I3(n24047), .O(n24049) );
  MUX2 U25534 ( .A(img[1871]), .B(n24049), .S(n28698), .O(n11661) );
  AOI22S U25535 ( .A1(n28106), .A2(img[1751]), .B1(n23941), .B2(n30073), .O(
        n24050) );
  ND2S U25536 ( .I1(n24340), .I2(n24050), .O(n24053) );
  NR2P U25537 ( .I1(n24051), .I2(n24111), .O(n24277) );
  NR2 U25538 ( .I1(n24692), .I2(n24277), .O(n24266) );
  ND2S U25539 ( .I1(n24266), .I2(n24758), .O(n24052) );
  AOI22S U25540 ( .A1(n27735), .A2(n30074), .B1(n24313), .B2(img[1711]), .O(
        n24055) );
  ND2S U25541 ( .I1(n13819), .I2(img[1775]), .O(n24054) );
  ND3S U25542 ( .I1(n24340), .I2(n24055), .I3(n24054), .O(n24056) );
  MUX2 U25543 ( .A(img[1751]), .B(n24056), .S(n28705), .O(n11781) );
  AOI22S U25544 ( .A1(n25810), .A2(img[1775]), .B1(n13781), .B2(n30075), .O(
        n24057) );
  ND2S U25545 ( .I1(n24340), .I2(n24057), .O(n24058) );
  AOI22S U25546 ( .A1(n29096), .A2(n30076), .B1(n24313), .B2(img[1687]), .O(
        n24060) );
  AOI22S U25547 ( .A1(n13770), .A2(img[1751]), .B1(img[1783]), .B2(n13782), 
        .O(n24059) );
  ND3S U25548 ( .I1(n24340), .I2(n24060), .I3(n24059), .O(n24061) );
  MUX2 U25549 ( .A(img[1775]), .B(n24061), .S(n28712), .O(n11763) );
  AOI22S U25550 ( .A1(n27957), .A2(img[1783]), .B1(n24374), .B2(n30077), .O(
        n24062) );
  ND2S U25551 ( .I1(n24340), .I2(n24062), .O(n24063) );
  AOI22S U25552 ( .A1(n28075), .A2(n30078), .B1(n24313), .B2(img[1679]), .O(
        n24065) );
  AOI22S U25553 ( .A1(n13905), .A2(img[1743]), .B1(img[1775]), .B2(n13782), 
        .O(n24064) );
  ND3S U25554 ( .I1(n24340), .I2(n24065), .I3(n24064), .O(n24066) );
  MUX2 U25555 ( .A(img[1783]), .B(n24066), .S(n28719), .O(n11749) );
  AOI22S U25556 ( .A1(n13780), .A2(img[1743]), .B1(n24374), .B2(n30079), .O(
        n24067) );
  ND2S U25557 ( .I1(n24340), .I2(n24067), .O(n24068) );
  MUX2 U25558 ( .A(n24068), .B(img[1719]), .S(n28722), .O(n11813) );
  AOI22S U25559 ( .A1(n25591), .A2(n30080), .B1(n28043), .B2(img[1719]), .O(
        n24070) );
  ND3S U25560 ( .I1(n24340), .I2(n24070), .I3(n24069), .O(n24071) );
  MUX2 U25561 ( .A(img[1743]), .B(n24071), .S(n28726), .O(n11795) );
  AOI22S U25562 ( .A1(n28840), .A2(img[1623]), .B1(n28862), .B2(n30081), .O(
        n24072) );
  ND2S U25563 ( .I1(n24340), .I2(n24072), .O(n24073) );
  MUX2 U25564 ( .A(n24073), .B(img[1583]), .S(n28729), .O(n11949) );
  AOI22S U25565 ( .A1(n28862), .A2(n30082), .B1(n28254), .B2(img[1583]), .O(
        n24075) );
  ND3S U25566 ( .I1(n24340), .I2(n24075), .I3(n24074), .O(n24076) );
  MUX2 U25567 ( .A(img[1623]), .B(n24076), .S(n28733), .O(n11915) );
  AOI22S U25568 ( .A1(n28106), .A2(img[1647]), .B1(n13781), .B2(n30083), .O(
        n24077) );
  ND2S U25569 ( .I1(n24340), .I2(n24077), .O(n24078) );
  MUX2 U25570 ( .A(n24078), .B(img[1559]), .S(n28736), .O(n11979) );
  AOI22S U25571 ( .A1(n25468), .A2(n30084), .B1(n24313), .B2(img[1559]), .O(
        n24080) );
  AOI22S U25572 ( .A1(n13899), .A2(img[1623]), .B1(img[1655]), .B2(n13782), 
        .O(n24079) );
  ND3S U25573 ( .I1(n24340), .I2(n24080), .I3(n24079), .O(n24082) );
  NR2 U25574 ( .I1(n24542), .I2(n24345), .O(n24081) );
  MUX2 U25575 ( .A(img[1647]), .B(n24082), .S(n28740), .O(n11885) );
  AOI22S U25576 ( .A1(n28442), .A2(img[1655]), .B1(n23941), .B2(n30085), .O(
        n24083) );
  ND2S U25577 ( .I1(n24340), .I2(n24083), .O(n24085) );
  NR2 U25578 ( .I1(n24726), .I2(n24304), .O(n24084) );
  AOI22S U25579 ( .A1(n29242), .A2(n30086), .B1(n26504), .B2(img[1551]), .O(
        n24087) );
  AOI22S U25580 ( .A1(n13899), .A2(img[1615]), .B1(img[1647]), .B2(n13782), 
        .O(n24086) );
  ND3S U25581 ( .I1(n24340), .I2(n24087), .I3(n24086), .O(n24089) );
  NR2 U25582 ( .I1(n24670), .I2(n24345), .O(n24088) );
  MUX2 U25583 ( .A(img[1655]), .B(n24089), .S(n28747), .O(n11883) );
  AOI22S U25584 ( .A1(n29072), .A2(img[1615]), .B1(n28695), .B2(n30087), .O(
        n24090) );
  ND2S U25585 ( .I1(n24340), .I2(n24090), .O(n24092) );
  MUX2 U25586 ( .A(n24092), .B(img[1591]), .S(n28750), .O(n11947) );
  AOI22S U25587 ( .A1(n28433), .A2(n30088), .B1(n24890), .B2(img[1591]), .O(
        n24094) );
  ND3S U25588 ( .I1(n24340), .I2(n24094), .I3(n24093), .O(n24095) );
  MUX2 U25589 ( .A(img[1615]), .B(n24095), .S(n28754), .O(n11917) );
  AOI22S U25590 ( .A1(n28840), .A2(img[1143]), .B1(n28614), .B2(n30089), .O(
        n24096) );
  ND2S U25591 ( .I1(n24340), .I2(n24096), .O(n24100) );
  AOI22S U25592 ( .A1(n24193), .A2(n30090), .B1(n24313), .B2(img[1039]), .O(
        n24102) );
  ND3S U25593 ( .I1(n24340), .I2(n24102), .I3(n24101), .O(n24103) );
  MUX2 U25594 ( .A(img[1143]), .B(n24103), .S(n28761), .O(n12395) );
  AOI22S U25595 ( .A1(n26855), .A2(img[1103]), .B1(n29530), .B2(n30091), .O(
        n24104) );
  ND2S U25596 ( .I1(n24340), .I2(n24104), .O(n24106) );
  MUX2 U25597 ( .A(n24106), .B(img[1079]), .S(n28764), .O(n12459) );
  AOI22S U25598 ( .A1(n13781), .A2(n30092), .B1(n24313), .B2(img[1079]), .O(
        n24108) );
  ND3S U25599 ( .I1(n24340), .I2(n24108), .I3(n24107), .O(n24109) );
  MUX2 U25600 ( .A(img[1103]), .B(n24109), .S(n28768), .O(n12429) );
  AOI22S U25601 ( .A1(n27990), .A2(img[2007]), .B1(n24374), .B2(n30093), .O(
        n24110) );
  ND2S U25602 ( .I1(n24340), .I2(n24110), .O(n24114) );
  NR2P U25603 ( .I1(n24112), .I2(n24111), .O(n24351) );
  NR2 U25604 ( .I1(n24692), .I2(n24351), .O(n24335) );
  ND2S U25605 ( .I1(n24335), .I2(n24758), .O(n24113) );
  AOI22S U25606 ( .A1(n25062), .A2(n30094), .B1(n28069), .B2(img[1967]), .O(
        n24116) );
  ND2S U25607 ( .I1(n13905), .I2(img[2031]), .O(n24115) );
  ND3S U25608 ( .I1(n24340), .I2(n24116), .I3(n24115), .O(n24117) );
  MUX2 U25609 ( .A(img[2007]), .B(n24117), .S(n28775), .O(n11525) );
  AOI22S U25610 ( .A1(n13780), .A2(img[2031]), .B1(n29397), .B2(n30095), .O(
        n24118) );
  ND2S U25611 ( .I1(n24340), .I2(n24118), .O(n24119) );
  MUX2 U25612 ( .A(n24119), .B(img[1943]), .S(n28778), .O(n11589) );
  AOI22S U25613 ( .A1(n28037), .A2(n30096), .B1(n26504), .B2(img[1943]), .O(
        n24121) );
  AOI22S U25614 ( .A1(n13904), .A2(img[2007]), .B1(img[2039]), .B2(n13782), 
        .O(n24120) );
  ND3S U25615 ( .I1(n24340), .I2(n24121), .I3(n24120), .O(n24122) );
  MUX2 U25616 ( .A(img[2031]), .B(n24122), .S(n28782), .O(n11507) );
  AOI22S U25617 ( .A1(n26970), .A2(img[2039]), .B1(n24193), .B2(n30097), .O(
        n24123) );
  ND2S U25618 ( .I1(n24340), .I2(n24123), .O(n24124) );
  MUX2 U25619 ( .A(img[1935]), .B(n24124), .S(n28785), .O(n11603) );
  AOI22S U25620 ( .A1(n29096), .A2(n30098), .B1(n28069), .B2(img[1935]), .O(
        n24126) );
  AOI22S U25621 ( .A1(n13903), .A2(img[1999]), .B1(img[2031]), .B2(n13782), 
        .O(n24125) );
  ND3S U25622 ( .I1(n24340), .I2(n24126), .I3(n24125), .O(n24127) );
  MUX2 U25623 ( .A(img[2039]), .B(n24127), .S(n28789), .O(n11493) );
  AOI22S U25624 ( .A1(n26101), .A2(img[1999]), .B1(n25062), .B2(n30099), .O(
        n24128) );
  ND2S U25625 ( .I1(n24340), .I2(n24128), .O(n24131) );
  ND2S U25626 ( .I1(n24335), .I2(n24748), .O(n24130) );
  AOI22S U25627 ( .A1(n28037), .A2(n30100), .B1(n28069), .B2(img[1975]), .O(
        n24133) );
  ND2S U25628 ( .I1(n13820), .I2(img[2039]), .O(n24132) );
  ND3S U25629 ( .I1(n24340), .I2(n24133), .I3(n24132), .O(n24135) );
  MUX2 U25630 ( .A(img[1999]), .B(n24135), .S(n28796), .O(n11539) );
  AOI22S U25631 ( .A1(n13777), .A2(img[543]), .B1(n24193), .B2(n30101), .O(
        n24136) );
  ND2S U25632 ( .I1(n24340), .I2(n24136), .O(n24137) );
  NR2 U25633 ( .I1(n24234), .I2(n24147), .O(n24346) );
  NR2 U25634 ( .I1(n24346), .I2(n24692), .O(n24213) );
  AO12 U25635 ( .B1(n24213), .B2(n24694), .A1(n24693), .O(n29286) );
  MUX2 U25636 ( .A(n24137), .B(img[615]), .S(n29286), .O(n12923) );
  AOI22S U25637 ( .A1(n28347), .A2(img[615]), .B1(n13781), .B2(n30102), .O(
        n24138) );
  ND2S U25638 ( .I1(n24340), .I2(n24138), .O(n24141) );
  NR2 U25639 ( .I1(n24640), .I2(n24669), .O(n24140) );
  NR2 U25640 ( .I1(n24233), .I2(n24139), .O(n24350) );
  AOI22S U25641 ( .A1(n27746), .A2(img[31]), .B1(n25591), .B2(n30103), .O(
        n24142) );
  ND2S U25642 ( .I1(n24340), .I2(n24142), .O(n24143) );
  MUX2 U25643 ( .A(img[103]), .B(n24143), .S(n29280), .O(n13435) );
  AOI22S U25644 ( .A1(n13780), .A2(img[103]), .B1(n29096), .B2(n30104), .O(
        n24144) );
  ND2S U25645 ( .I1(n24340), .I2(n24144), .O(n24145) );
  NR2 U25646 ( .I1(n24350), .I2(n24692), .O(n24184) );
  AOI22S U25647 ( .A1(n28442), .A2(img[1247]), .B1(n27443), .B2(n30105), .O(
        n24146) );
  ND2S U25648 ( .I1(n24340), .I2(n24146), .O(n24149) );
  NR2 U25649 ( .I1(n24147), .I2(n24220), .O(n24619) );
  NR2 U25650 ( .I1(n24619), .I2(n24692), .O(n24612) );
  MUX2 U25651 ( .A(n24149), .B(img[1191]), .S(n29207), .O(n12341) );
  AOI22S U25652 ( .A1(n13779), .A2(n30106), .B1(n25444), .B2(img[1191]), .O(
        n24151) );
  ND3S U25653 ( .I1(n24340), .I2(n24151), .I3(n24150), .O(n24154) );
  INV1S U25654 ( .I(n24152), .O(n24153) );
  NR2 U25655 ( .I1(n24233), .I2(n24153), .O(n24622) );
  MUX2 U25656 ( .A(img[1247]), .B(n24154), .S(n29211), .O(n12291) );
  AOI22S U25657 ( .A1(n29194), .A2(n30107), .B1(n28069), .B2(img[1183]), .O(
        n24156) );
  ND3S U25658 ( .I1(n24340), .I2(n24156), .I3(n24155), .O(n24157) );
  MUX2 U25659 ( .A(img[1255]), .B(n24157), .S(n29218), .O(n12277) );
  AOI22S U25660 ( .A1(n29072), .A2(img[1255]), .B1(n28862), .B2(n30108), .O(
        n24158) );
  ND2S U25661 ( .I1(n24340), .I2(n24158), .O(n24160) );
  NR2 U25662 ( .I1(n24463), .I2(n24669), .O(n24159) );
  AOI22S U25663 ( .A1(n28347), .A2(img[1375]), .B1(n29457), .B2(n30109), .O(
        n24161) );
  ND2S U25664 ( .I1(n24340), .I2(n24161), .O(n24162) );
  MUX2 U25665 ( .A(n24162), .B(img[1319]), .S(n29233), .O(n12219) );
  AOI22S U25666 ( .A1(n29096), .A2(n30110), .B1(n28254), .B2(img[1319]), .O(
        n24164) );
  ND2S U25667 ( .I1(n29124), .I2(img[1383]), .O(n24163) );
  ND3S U25668 ( .I1(n24340), .I2(n24164), .I3(n24163), .O(n24165) );
  MUX2 U25669 ( .A(img[1375]), .B(n24165), .S(n29237), .O(n12157) );
  AOI22S U25670 ( .A1(n29096), .A2(n30111), .B1(n28069), .B2(img[1311]), .O(
        n24167) );
  ND3S U25671 ( .I1(n24340), .I2(n24167), .I3(n24166), .O(n24168) );
  MUX2 U25672 ( .A(img[1383]), .B(n24168), .S(n29245), .O(n12155) );
  AOI22S U25673 ( .A1(n27990), .A2(img[1383]), .B1(n28614), .B2(n30112), .O(
        n24169) );
  ND2S U25674 ( .I1(n24340), .I2(n24169), .O(n24170) );
  MUX2 U25675 ( .A(img[1311]), .B(n24170), .S(n29240), .O(n12221) );
  AOI22S U25676 ( .A1(n27990), .A2(img[927]), .B1(n29242), .B2(n30113), .O(
        n24171) );
  ND2S U25677 ( .I1(n24340), .I2(n24171), .O(n24173) );
  NR2 U25678 ( .I1(n24346), .I2(n24716), .O(n24172) );
  NR2P U25679 ( .I1(n24172), .I2(n24717), .O(n29224) );
  MUX2 U25680 ( .A(img[999]), .B(n24173), .S(n29224), .O(n12533) );
  AOI22S U25681 ( .A1(n13778), .A2(img[999]), .B1(n24755), .B2(n30114), .O(
        n24174) );
  ND2S U25682 ( .I1(n24340), .I2(n24174), .O(n24176) );
  NR2 U25683 ( .I1(n24646), .I2(n24669), .O(n24175) );
  AOI22S U25684 ( .A1(n28382), .A2(img[159]), .B1(n23941), .B2(n30115), .O(
        n24177) );
  ND2S U25685 ( .I1(n24340), .I2(n24177), .O(n24178) );
  MUX2 U25686 ( .A(img[231]), .B(n24178), .S(n29267), .O(n13301) );
  AOI22S U25687 ( .A1(n26855), .A2(img[231]), .B1(n23941), .B2(n30116), .O(
        n24179) );
  ND2S U25688 ( .I1(n24340), .I2(n24179), .O(n24180) );
  MUX2 U25689 ( .A(img[159]), .B(n24180), .S(n29264), .O(n13379) );
  AOI22S U25690 ( .A1(n28083), .A2(img[287]), .B1(n23941), .B2(n30117), .O(
        n24181) );
  ND2S U25691 ( .I1(n24340), .I2(n24181), .O(n24182) );
  OAI12HS U25692 ( .B1(n24732), .B2(n24213), .A1(n24495), .O(n29182) );
  MUX2 U25693 ( .A(img[359]), .B(n24182), .S(n29182), .O(n13179) );
  AOI22S U25694 ( .A1(n29072), .A2(img[359]), .B1(n23941), .B2(n30118), .O(
        n24183) );
  ND2S U25695 ( .I1(n24340), .I2(n24183), .O(n24185) );
  OAI12HS U25696 ( .B1(n24732), .B2(n24184), .A1(n24495), .O(n29179) );
  BUF2 U25697 ( .I(n24581), .O(n24349) );
  AOI22S U25698 ( .A1(n28840), .A2(img[415]), .B1(n23941), .B2(n30119), .O(
        n24186) );
  ND2S U25699 ( .I1(n24349), .I2(n24186), .O(n24187) );
  MUX2 U25700 ( .A(img[487]), .B(n24187), .S(n29273), .O(n13045) );
  AOI22S U25701 ( .A1(n13773), .A2(img[487]), .B1(n23941), .B2(n30120), .O(
        n24188) );
  ND2S U25702 ( .I1(n24349), .I2(n24188), .O(n24189) );
  NR2P U25703 ( .I1(n24319), .I2(n24740), .O(n29270) );
  MUX2 U25704 ( .A(img[415]), .B(n24189), .S(n29270), .O(n13123) );
  AOI22S U25705 ( .A1(n26822), .A2(img[1503]), .B1(n23941), .B2(n30121), .O(
        n24190) );
  ND2S U25706 ( .I1(n24349), .I2(n24190), .O(n24192) );
  ND2S U25707 ( .I1(n24520), .I2(n24694), .O(n24191) );
  ND2 U25708 ( .I1(n24633), .I2(n24191), .O(n29248) );
  MUX2 U25709 ( .A(n24192), .B(img[1447]), .S(n29248), .O(n12085) );
  AOI22S U25710 ( .A1(n29194), .A2(n30122), .B1(n25444), .B2(img[1447]), .O(
        n24195) );
  ND3S U25711 ( .I1(n24340), .I2(n24195), .I3(n24194), .O(n24197) );
  AOI22S U25712 ( .A1(n29194), .A2(n30123), .B1(n24313), .B2(img[1439]), .O(
        n24199) );
  ND2S U25713 ( .I1(n13770), .I2(img[1503]), .O(n24198) );
  ND3S U25714 ( .I1(n24340), .I2(n24199), .I3(n24198), .O(n24201) );
  MUX2 U25715 ( .A(img[1511]), .B(n24201), .S(n29261), .O(n12021) );
  AOI22S U25716 ( .A1(n28382), .A2(img[1511]), .B1(n23941), .B2(n30124), .O(
        n24202) );
  ND2S U25717 ( .I1(n24349), .I2(n24202), .O(n24204) );
  MUX2 U25718 ( .A(n24204), .B(img[1439]), .S(n29255), .O(n12099) );
  INV1S U25719 ( .I(img[871]), .O(n24205) );
  AOI22S U25720 ( .A1(n13773), .A2(img[799]), .B1(n29096), .B2(n24205), .O(
        n24206) );
  ND2S U25721 ( .I1(n24349), .I2(n24206), .O(n24208) );
  ND2S U25722 ( .I1(n24748), .I2(n24213), .O(n24207) );
  AOI22S U25723 ( .A1(n26822), .A2(img[871]), .B1(n13781), .B2(n30125), .O(
        n24209) );
  ND2S U25724 ( .I1(n24349), .I2(n24209), .O(n24211) );
  NR2 U25725 ( .I1(n24673), .I2(n24669), .O(n24210) );
  MUX2 U25726 ( .A(img[799]), .B(n24211), .S(n29227), .O(n12733) );
  AOI22S U25727 ( .A1(n13773), .A2(img[671]), .B1(n13775), .B2(n30126), .O(
        n24212) );
  ND2S U25728 ( .I1(n24349), .I2(n24212), .O(n24215) );
  ND2S U25729 ( .I1(n24758), .I2(n24213), .O(n24214) );
  AOI22S U25730 ( .A1(n28382), .A2(img[743]), .B1(n28862), .B2(n30127), .O(
        n24216) );
  ND2S U25731 ( .I1(n24349), .I2(n24216), .O(n24218) );
  NR2 U25732 ( .I1(n24681), .I2(n24669), .O(n24217) );
  MUX2 U25733 ( .A(img[671]), .B(n24218), .S(n29201), .O(n12867) );
  AOI22S U25734 ( .A1(n27746), .A2(img[1863]), .B1(n29242), .B2(n30128), .O(
        n24219) );
  ND2S U25735 ( .I1(n24349), .I2(n24219), .O(n24221) );
  NR2 U25736 ( .I1(n24233), .I2(n24220), .O(n24398) );
  MUX2 U25737 ( .A(img[1855]), .B(n24221), .S(n28919), .O(n11677) );
  AOI22S U25738 ( .A1(n25062), .A2(n30129), .B1(n28069), .B2(img[1855]), .O(
        n24223) );
  ND2S U25739 ( .I1(n13770), .I2(img[1919]), .O(n24222) );
  ND3S U25740 ( .I1(n24340), .I2(n24223), .I3(n24222), .O(n24224) );
  MUX2 U25741 ( .A(img[1863]), .B(n24224), .S(n28916), .O(n11675) );
  AOI22S U25742 ( .A1(n13777), .A2(img[1919]), .B1(n13781), .B2(n30130), .O(
        n24225) );
  ND2S U25743 ( .I1(n24349), .I2(n24225), .O(n24230) );
  INV1S U25744 ( .I(n24226), .O(n24227) );
  NR2 U25745 ( .I1(n24228), .I2(n24227), .O(n24708) );
  AOI22S U25746 ( .A1(n25062), .A2(n30131), .B1(n28069), .B2(img[1799]), .O(
        n24232) );
  AOI22S U25747 ( .A1(n13899), .A2(img[1863]), .B1(img[1895]), .B2(n13782), 
        .O(n24231) );
  ND3S U25748 ( .I1(n24340), .I2(n24232), .I3(n24231), .O(n24236) );
  NR2 U25749 ( .I1(n24234), .I2(n24233), .O(n24727) );
  MUX2 U25750 ( .A(img[1919]), .B(n24236), .S(n28911), .O(n11613) );
  AOI22S U25751 ( .A1(n28083), .A2(img[1887]), .B1(n28862), .B2(n30132), .O(
        n24237) );
  ND2S U25752 ( .I1(n24349), .I2(n24237), .O(n24241) );
  NR2 U25753 ( .I1(n24612), .I2(n24238), .O(n24239) );
  NR2 U25754 ( .I1(n24240), .I2(n24239), .O(n28892) );
  MUX2 U25755 ( .A(n24241), .B(img[1831]), .S(n28892), .O(n11707) );
  AOI22S U25756 ( .A1(n28075), .A2(n30133), .B1(n27919), .B2(img[1831]), .O(
        n24243) );
  ND3S U25757 ( .I1(n24340), .I2(n24243), .I3(n24242), .O(n24245) );
  AOI22S U25758 ( .A1(n28135), .A2(n30134), .B1(n24313), .B2(img[1823]), .O(
        n24247) );
  AOI22S U25759 ( .A1(n13903), .A2(img[1887]), .B1(img[1919]), .B2(n13782), 
        .O(n24246) );
  ND3S U25760 ( .I1(n24340), .I2(n24247), .I3(n24246), .O(n24248) );
  MUX2 U25761 ( .A(img[1895]), .B(n24248), .S(n28903), .O(n11643) );
  AOI22S U25762 ( .A1(n27990), .A2(img[1895]), .B1(n29397), .B2(n30135), .O(
        n24249) );
  ND2S U25763 ( .I1(n24349), .I2(n24249), .O(n24252) );
  NR2 U25764 ( .I1(n24669), .I2(n24250), .O(n24251) );
  MUX2 U25765 ( .A(img[1823]), .B(n24252), .S(n28899), .O(n11709) );
  AOI22S U25766 ( .A1(n28347), .A2(img[1735]), .B1(n28433), .B2(n30136), .O(
        n24253) );
  ND2S U25767 ( .I1(n24349), .I2(n24253), .O(n24255) );
  NR2 U25768 ( .I1(n24398), .I2(n24716), .O(n24440) );
  NR2 U25769 ( .I1(n24716), .I2(n24277), .O(n24254) );
  MUX2 U25770 ( .A(img[1727]), .B(n24255), .S(n28948), .O(n11811) );
  AOI22S U25771 ( .A1(n29242), .A2(n30137), .B1(n24313), .B2(img[1727]), .O(
        n24257) );
  ND3S U25772 ( .I1(n24340), .I2(n24257), .I3(n24256), .O(n24258) );
  MUX2 U25773 ( .A(img[1735]), .B(n24258), .S(n28945), .O(n11797) );
  AOI22S U25774 ( .A1(n26822), .A2(img[1791]), .B1(n25859), .B2(n30138), .O(
        n24259) );
  ND2S U25775 ( .I1(n24349), .I2(n24259), .O(n24260) );
  AOI22S U25776 ( .A1(n23941), .A2(n30139), .B1(n24313), .B2(img[1671]), .O(
        n24262) );
  AOI22S U25777 ( .A1(n13903), .A2(img[1735]), .B1(img[1767]), .B2(n13782), 
        .O(n24261) );
  ND3S U25778 ( .I1(n24340), .I2(n24262), .I3(n24261), .O(n24264) );
  MUX2 U25779 ( .A(img[1791]), .B(n24264), .S(n28941), .O(n11747) );
  AOI22S U25780 ( .A1(n29129), .A2(img[1759]), .B1(n28862), .B2(n30140), .O(
        n24265) );
  ND2S U25781 ( .I1(n24349), .I2(n24265), .O(n24268) );
  ND2S U25782 ( .I1(n24266), .I2(n24694), .O(n24267) );
  MUX2 U25783 ( .A(n24268), .B(img[1703]), .S(n28922), .O(n11829) );
  AOI22S U25784 ( .A1(n24374), .A2(n30141), .B1(n24313), .B2(img[1703]), .O(
        n24270) );
  ND3S U25785 ( .I1(n24340), .I2(n24270), .I3(n24269), .O(n24272) );
  AOI22S U25786 ( .A1(n13781), .A2(n30142), .B1(n24313), .B2(img[1695]), .O(
        n24274) );
  AOI22S U25787 ( .A1(n13904), .A2(img[1759]), .B1(img[1791]), .B2(n13782), 
        .O(n24273) );
  ND3S U25788 ( .I1(n24340), .I2(n24274), .I3(n24273), .O(n24275) );
  MUX2 U25789 ( .A(img[1767]), .B(n24275), .S(n28933), .O(n11765) );
  AOI22S U25790 ( .A1(n13777), .A2(img[1767]), .B1(n28862), .B2(n30143), .O(
        n24276) );
  ND2S U25791 ( .I1(n24349), .I2(n24276), .O(n24278) );
  MUX2 U25792 ( .A(img[1695]), .B(n24278), .S(n28929), .O(n11843) );
  AOI22S U25793 ( .A1(n13777), .A2(img[1607]), .B1(n25591), .B2(n30144), .O(
        n24279) );
  ND2S U25794 ( .I1(n24349), .I2(n24279), .O(n24281) );
  NR2 U25795 ( .I1(n24716), .I2(n24304), .O(n24280) );
  AOI22S U25796 ( .A1(n29397), .A2(n30145), .B1(n24313), .B2(img[1599]), .O(
        n24283) );
  ND2S U25797 ( .I1(n13820), .I2(img[1663]), .O(n24282) );
  ND3S U25798 ( .I1(n24340), .I2(n24283), .I3(n24282), .O(n24284) );
  MUX2 U25799 ( .A(img[1607]), .B(n24284), .S(n28973), .O(n11931) );
  AOI22S U25800 ( .A1(n28106), .A2(img[1663]), .B1(n25062), .B2(n30146), .O(
        n24285) );
  ND2S U25801 ( .I1(n24349), .I2(n24285), .O(n24286) );
  AOI22S U25802 ( .A1(n29194), .A2(n30147), .B1(n24313), .B2(img[1543]), .O(
        n24288) );
  AOI22S U25803 ( .A1(n13899), .A2(img[1607]), .B1(img[1639]), .B2(n13782), 
        .O(n24287) );
  ND3S U25804 ( .I1(n24340), .I2(n24288), .I3(n24287), .O(n24291) );
  NR2 U25805 ( .I1(n24727), .I2(n24345), .O(n24290) );
  MUX2 U25806 ( .A(img[1663]), .B(n24291), .S(n28969), .O(n11869) );
  AOI22S U25807 ( .A1(n27990), .A2(img[1631]), .B1(n13781), .B2(n30148), .O(
        n24292) );
  ND2S U25808 ( .I1(n24349), .I2(n24292), .O(n24295) );
  MUX2 U25809 ( .A(n24295), .B(img[1575]), .S(n28951), .O(n11963) );
  AOI22S U25810 ( .A1(n28695), .A2(n30149), .B1(n24313), .B2(img[1575]), .O(
        n24297) );
  ND2S U25811 ( .I1(n13770), .I2(img[1639]), .O(n24296) );
  ND3S U25812 ( .I1(n24340), .I2(n24297), .I3(n24296), .O(n24299) );
  AOI22S U25813 ( .A1(n28938), .A2(n30150), .B1(n24313), .B2(img[1567]), .O(
        n24301) );
  AOI22S U25814 ( .A1(n29124), .A2(img[1631]), .B1(img[1663]), .B2(n13782), 
        .O(n24300) );
  ND3S U25815 ( .I1(n24340), .I2(n24301), .I3(n24300), .O(n24302) );
  MUX2 U25816 ( .A(img[1639]), .B(n24302), .S(n28962), .O(n11898) );
  AOI22S U25817 ( .A1(n29072), .A2(img[1639]), .B1(n28135), .B2(n30151), .O(
        n24303) );
  ND2S U25818 ( .I1(n24349), .I2(n24303), .O(n24306) );
  NR2 U25819 ( .I1(n24669), .I2(n24304), .O(n24305) );
  MUX2 U25820 ( .A(img[1567]), .B(n24306), .S(n28958), .O(n11965) );
  AOI22S U25821 ( .A1(n28347), .A2(img[1119]), .B1(n28862), .B2(n30152), .O(
        n24307) );
  ND2S U25822 ( .I1(n24349), .I2(n24307), .O(n24309) );
  MUX2 U25823 ( .A(n24309), .B(img[1063]), .S(n29185), .O(n12475) );
  AOI22S U25824 ( .A1(n29194), .A2(n30153), .B1(n24313), .B2(img[1063]), .O(
        n24311) );
  ND3S U25825 ( .I1(n24340), .I2(n24311), .I3(n24310), .O(n24312) );
  MUX2 U25826 ( .A(img[1119]), .B(n24312), .S(n29189), .O(n12413) );
  AOI22S U25827 ( .A1(n28162), .A2(n30154), .B1(n24313), .B2(img[1055]), .O(
        n24315) );
  ND2S U25828 ( .I1(n13770), .I2(img[1119]), .O(n24314) );
  ND3S U25829 ( .I1(n24340), .I2(n24315), .I3(n24314), .O(n24316) );
  MUX2 U25830 ( .A(img[1127]), .B(n24316), .S(n29198), .O(n12411) );
  AOI22S U25831 ( .A1(n13771), .A2(img[1127]), .B1(n13781), .B2(n30155), .O(
        n24317) );
  ND2S U25832 ( .I1(n24349), .I2(n24317), .O(n24320) );
  NR2 U25833 ( .I1(n24669), .I2(n24543), .O(n24318) );
  AOI22S U25834 ( .A1(n29435), .A2(img[1991]), .B1(n13781), .B2(n30156), .O(
        n24321) );
  ND2S U25835 ( .I1(n24349), .I2(n24321), .O(n24322) );
  MUX2 U25836 ( .A(img[1983]), .B(n24322), .S(n29018), .O(n11555) );
  AOI22S U25837 ( .A1(n27735), .A2(n30157), .B1(n24434), .B2(img[1983]), .O(
        n24324) );
  ND2S U25838 ( .I1(n29124), .I2(img[2047]), .O(n24323) );
  ND3 U25839 ( .I1(n24581), .I2(n24324), .I3(n24323), .O(n24325) );
  AOI22S U25840 ( .A1(n24415), .A2(img[2047]), .B1(n24755), .B2(n30158), .O(
        n24326) );
  ND2S U25841 ( .I1(n24349), .I2(n24326), .O(n24327) );
  MUX2 U25842 ( .A(img[1927]), .B(n24327), .S(n29007), .O(n11605) );
  AOI22S U25843 ( .A1(n25062), .A2(n30159), .B1(n24434), .B2(img[1927]), .O(
        n24329) );
  AOI22S U25844 ( .A1(n13904), .A2(img[1991]), .B1(img[2023]), .B2(n13782), 
        .O(n24328) );
  INV1S U25845 ( .I(n24345), .O(n24330) );
  OAI112HS U25846 ( .C1(n24332), .C2(n24699), .A1(n24331), .B1(n24330), .O(
        n29011) );
  AOI22S U25847 ( .A1(n24415), .A2(img[2015]), .B1(n29530), .B2(n30160), .O(
        n24334) );
  ND2S U25848 ( .I1(n24349), .I2(n24334), .O(n24337) );
  ND2S U25849 ( .I1(n24335), .I2(n24694), .O(n24336) );
  MUX2 U25850 ( .A(n24337), .B(img[1959]), .S(n28993), .O(n11573) );
  AOI22S U25851 ( .A1(n27443), .A2(n30161), .B1(n24434), .B2(img[1959]), .O(
        n24339) );
  ND3S U25852 ( .I1(n24340), .I2(n24339), .I3(n24338), .O(n24342) );
  AOI22S U25853 ( .A1(n29194), .A2(n30162), .B1(n24434), .B2(img[1951]), .O(
        n24344) );
  AOI22S U25854 ( .A1(n13770), .A2(img[2015]), .B1(img[2047]), .B2(n13782), 
        .O(n24343) );
  ND3S U25855 ( .I1(n24340), .I2(n24344), .I3(n24343), .O(n24347) );
  MUX2 U25856 ( .A(img[2023]), .B(n24347), .S(n29004), .O(n11509) );
  AOI22S U25857 ( .A1(n24415), .A2(img[2023]), .B1(n24755), .B2(n30163), .O(
        n24348) );
  ND2S U25858 ( .I1(n24349), .I2(n24348), .O(n24352) );
  MUX2 U25859 ( .A(img[1951]), .B(n24352), .S(n29000), .O(n11587) );
  BUF2 U25860 ( .I(n24581), .O(n24424) );
  AOI22S U25861 ( .A1(n24415), .A2(img[583]), .B1(n25062), .B2(n30164), .O(
        n24353) );
  ND2S U25862 ( .I1(n24424), .I2(n24353), .O(n24354) );
  NR2 U25863 ( .I1(n24398), .I2(n24692), .O(n24425) );
  AO12 U25864 ( .B1(n24425), .B2(n24694), .A1(n24693), .O(n29532) );
  MUX2 U25865 ( .A(n24354), .B(img[575]), .S(n29532), .O(n12957) );
  AOI22S U25866 ( .A1(n28347), .A2(img[575]), .B1(n28695), .B2(n30165), .O(
        n24355) );
  ND2S U25867 ( .I1(n24424), .I2(n24355), .O(n24356) );
  NR2 U25868 ( .I1(n24444), .I2(n24692), .O(n24429) );
  AO12 U25869 ( .B1(n24429), .B2(n24694), .A1(n24693), .O(n28799) );
  MUX2 U25870 ( .A(n24356), .B(img[583]), .S(n28799), .O(n12955) );
  AOI22S U25871 ( .A1(n28840), .A2(img[71]), .B1(n28182), .B2(n30166), .O(
        n24357) );
  ND2S U25872 ( .I1(n24424), .I2(n24357), .O(n24358) );
  AOI22S U25873 ( .A1(n13778), .A2(img[63]), .B1(n28938), .B2(n30167), .O(
        n24359) );
  ND2S U25874 ( .I1(n24424), .I2(n24359), .O(n24360) );
  MUX2 U25875 ( .A(img[71]), .B(n24360), .S(n28804), .O(n13467) );
  AOI22S U25876 ( .A1(n28347), .A2(img[1279]), .B1(n29530), .B2(n30168), .O(
        n24361) );
  ND2S U25877 ( .I1(n24424), .I2(n24361), .O(n24362) );
  NR2P U25878 ( .I1(n24229), .I2(n24466), .O(n28810) );
  MUX2 U25879 ( .A(img[1159]), .B(n24362), .S(n28810), .O(n12373) );
  AOI22S U25880 ( .A1(n29194), .A2(n30169), .B1(n24434), .B2(img[1159]), .O(
        n24364) );
  ND3S U25881 ( .I1(n24340), .I2(n24364), .I3(n24363), .O(n24365) );
  MUX2 U25882 ( .A(img[1279]), .B(n24365), .S(n28814), .O(n12259) );
  AOI22S U25883 ( .A1(n25595), .A2(img[1223]), .B1(n28075), .B2(n30170), .O(
        n24366) );
  ND2S U25884 ( .I1(n24424), .I2(n24366), .O(n24368) );
  MUX2 U25885 ( .A(img[1215]), .B(n24368), .S(n28821), .O(n12323) );
  AOI22S U25886 ( .A1(n29194), .A2(n30171), .B1(n24434), .B2(img[1215]), .O(
        n24370) );
  ND2S U25887 ( .I1(n13819), .I2(img[1279]), .O(n24369) );
  ND3S U25888 ( .I1(n24340), .I2(n24370), .I3(n24369), .O(n24371) );
  MUX2 U25889 ( .A(img[1223]), .B(n24371), .S(n28818), .O(n12309) );
  AOI22S U25890 ( .A1(n13772), .A2(img[1407]), .B1(n29457), .B2(n30172), .O(
        n24372) );
  ND2S U25891 ( .I1(n24424), .I2(n24372), .O(n24373) );
  AOI22S U25892 ( .A1(n28614), .A2(n30173), .B1(n24434), .B2(img[1287]), .O(
        n24376) );
  ND2S U25893 ( .I1(n13770), .I2(img[1351]), .O(n24375) );
  ND3S U25894 ( .I1(n24340), .I2(n24376), .I3(n24375), .O(n24377) );
  MUX2 U25895 ( .A(img[1407]), .B(n24377), .S(n28828), .O(n12125) );
  AOI22S U25896 ( .A1(n28382), .A2(img[1351]), .B1(n29242), .B2(n30174), .O(
        n24378) );
  ND2S U25897 ( .I1(n24424), .I2(n24378), .O(n24380) );
  NR2 U25898 ( .I1(n24716), .I2(n24476), .O(n24379) );
  MUX2 U25899 ( .A(img[1343]), .B(n24380), .S(n28835), .O(n12189) );
  AOI22S U25900 ( .A1(n28343), .A2(n30175), .B1(n24434), .B2(img[1343]), .O(
        n24382) );
  ND3S U25901 ( .I1(n24340), .I2(n24382), .I3(n24381), .O(n24383) );
  MUX2 U25902 ( .A(img[1351]), .B(n24383), .S(n28832), .O(n12187) );
  AOI22S U25903 ( .A1(n27746), .A2(img[967]), .B1(n28913), .B2(n30176), .O(
        n24384) );
  ND2S U25904 ( .I1(n24424), .I2(n24384), .O(n24385) );
  NR2P U25905 ( .I1(n24717), .I2(n24440), .O(n28842) );
  MUX2 U25906 ( .A(img[959]), .B(n24385), .S(n28842), .O(n12579) );
  AOI22S U25907 ( .A1(n28442), .A2(img[959]), .B1(n24755), .B2(n30177), .O(
        n24386) );
  ND2S U25908 ( .I1(n24424), .I2(n24386), .O(n24388) );
  NR2 U25909 ( .I1(n24444), .I2(n24716), .O(n24387) );
  NR2P U25910 ( .I1(n24387), .I2(n24717), .O(n28838) );
  AOI22S U25911 ( .A1(n29414), .A2(img[199]), .B1(n13779), .B2(n30178), .O(
        n24389) );
  ND2S U25912 ( .I1(n24424), .I2(n24389), .O(n24390) );
  MUX2 U25913 ( .A(img[191]), .B(n24390), .S(n28848), .O(n13347) );
  AOI22S U25914 ( .A1(n26822), .A2(img[191]), .B1(n24755), .B2(n30179), .O(
        n24391) );
  ND2S U25915 ( .I1(n24424), .I2(n24391), .O(n24392) );
  MUX2 U25916 ( .A(img[199]), .B(n24392), .S(n28845), .O(n13333) );
  AOI22S U25917 ( .A1(n24415), .A2(img[327]), .B1(n13781), .B2(n30180), .O(
        n24393) );
  ND2S U25918 ( .I1(n24424), .I2(n24393), .O(n24394) );
  OAI12HS U25919 ( .B1(n24732), .B2(n24425), .A1(n24495), .O(n28854) );
  AOI22S U25920 ( .A1(n24415), .A2(img[319]), .B1(n28695), .B2(n30181), .O(
        n24395) );
  ND2S U25921 ( .I1(n24424), .I2(n24395), .O(n24396) );
  OAI12HS U25922 ( .B1(n24732), .B2(n24429), .A1(n24495), .O(n28851) );
  MUX2 U25923 ( .A(img[327]), .B(n24396), .S(n28851), .O(n13211) );
  AOI22S U25924 ( .A1(n24415), .A2(img[455]), .B1(n27735), .B2(n30182), .O(
        n24397) );
  ND2S U25925 ( .I1(n24424), .I2(n24397), .O(n24399) );
  OA12 U25926 ( .B1(n24398), .B2(n24669), .A1(n24668), .O(n28860) );
  AOI22S U25927 ( .A1(n24415), .A2(img[447]), .B1(n23941), .B2(n30183), .O(
        n24400) );
  ND2S U25928 ( .I1(n24424), .I2(n24400), .O(n24401) );
  MUX2 U25929 ( .A(img[455]), .B(n24401), .S(n28857), .O(n13077) );
  AOI22S U25930 ( .A1(n24415), .A2(img[1535]), .B1(n13781), .B2(n30184), .O(
        n24402) );
  ND2S U25931 ( .I1(n24424), .I2(n24402), .O(n24403) );
  AOI22S U25932 ( .A1(n28343), .A2(n30185), .B1(n24434), .B2(img[1415]), .O(
        n24405) );
  ND2S U25933 ( .I1(n13770), .I2(img[1479]), .O(n24404) );
  ND3S U25934 ( .I1(n24340), .I2(n24405), .I3(n24404), .O(n24407) );
  MUX2 U25935 ( .A(img[1535]), .B(n24407), .S(n28868), .O(n12003) );
  AOI22S U25936 ( .A1(n24415), .A2(img[1479]), .B1(n25062), .B2(n30186), .O(
        n24408) );
  ND2S U25937 ( .I1(n24424), .I2(n24408), .O(n24410) );
  NR2 U25938 ( .I1(n24515), .I2(n24716), .O(n24409) );
  AOI22S U25939 ( .A1(n28037), .A2(n30187), .B1(n24434), .B2(img[1471]), .O(
        n24412) );
  ND2S U25940 ( .I1(n13770), .I2(img[1535]), .O(n24411) );
  ND3S U25941 ( .I1(n24340), .I2(n24412), .I3(n24411), .O(n24413) );
  MUX2 U25942 ( .A(img[1479]), .B(n24413), .S(n28872), .O(n12053) );
  INV1S U25943 ( .I(img[831]), .O(n24414) );
  AOI22S U25944 ( .A1(n24415), .A2(img[839]), .B1(n23941), .B2(n24414), .O(
        n24416) );
  ND2S U25945 ( .I1(n24424), .I2(n24416), .O(n24418) );
  ND2S U25946 ( .I1(n24748), .I2(n24425), .O(n24417) );
  INV1S U25947 ( .I(img[839]), .O(n24419) );
  AOI22S U25948 ( .A1(n27065), .A2(img[831]), .B1(n23918), .B2(n24419), .O(
        n24420) );
  ND2S U25949 ( .I1(n24424), .I2(n24420), .O(n24422) );
  ND2S U25950 ( .I1(n24748), .I2(n24429), .O(n24421) );
  MUX2 U25951 ( .A(n24422), .B(img[839]), .S(n28879), .O(n12699) );
  AOI22S U25952 ( .A1(n29072), .A2(img[711]), .B1(n28862), .B2(n30188), .O(
        n24423) );
  ND2S U25953 ( .I1(n24424), .I2(n24423), .O(n24427) );
  ND2S U25954 ( .I1(n24758), .I2(n24425), .O(n24426) );
  AOI22S U25955 ( .A1(n24415), .A2(img[703]), .B1(n23941), .B2(n30189), .O(
        n24428) );
  ND2S U25956 ( .I1(n24340), .I2(n24428), .O(n24431) );
  ND2S U25957 ( .I1(n24758), .I2(n24429), .O(n24430) );
  AOI22S U25958 ( .A1(n28347), .A2(img[1151]), .B1(n23941), .B2(n30190), .O(
        n24432) );
  ND2S U25959 ( .I1(n24340), .I2(n24432), .O(n24433) );
  MUX2 U25960 ( .A(img[1031]), .B(n24433), .S(n28979), .O(n12507) );
  AOI22S U25961 ( .A1(n13779), .A2(n30191), .B1(n24434), .B2(img[1031]), .O(
        n24436) );
  ND3S U25962 ( .I1(n24340), .I2(n24436), .I3(n24435), .O(n24437) );
  MUX2 U25963 ( .A(img[1151]), .B(n24437), .S(n28983), .O(n12381) );
  AOI22S U25964 ( .A1(n26101), .A2(img[1095]), .B1(n25062), .B2(n30192), .O(
        n24438) );
  ND2S U25965 ( .I1(n24340), .I2(n24438), .O(n24441) );
  NR2 U25966 ( .I1(n24716), .I2(n24543), .O(n24439) );
  AOI22S U25967 ( .A1(n13779), .A2(n30193), .B1(n24808), .B2(img[1087]), .O(
        n24443) );
  ND2S U25968 ( .I1(n13770), .I2(img[1151]), .O(n24442) );
  ND3S U25969 ( .I1(n24340), .I2(n24443), .I3(n24442), .O(n24445) );
  MUX2 U25970 ( .A(img[1095]), .B(n24445), .S(n28987), .O(n12440) );
  AOI22S U25971 ( .A1(n28318), .A2(img[535]), .B1(n24374), .B2(n30194), .O(
        n24446) );
  ND2S U25972 ( .I1(n24424), .I2(n24446), .O(n24447) );
  NR2 U25973 ( .I1(n24542), .I2(n24692), .O(n24529) );
  AO12 U25974 ( .B1(n24529), .B2(n24694), .A1(n24693), .O(n29024) );
  MUX2 U25975 ( .A(n24447), .B(img[623]), .S(n29024), .O(n12909) );
  AOI22S U25976 ( .A1(n27746), .A2(img[623]), .B1(n28862), .B2(n30195), .O(
        n24448) );
  ND2S U25977 ( .I1(n24340), .I2(n24448), .O(n24450) );
  INV1S U25978 ( .I(n24023), .O(n24500) );
  AOI22S U25979 ( .A1(n25810), .A2(img[23]), .B1(n25377), .B2(n30196), .O(
        n24451) );
  ND2S U25980 ( .I1(n24424), .I2(n24451), .O(n24452) );
  MUX2 U25981 ( .A(img[111]), .B(n24452), .S(n29030), .O(n13421) );
  AOI22S U25982 ( .A1(n28347), .A2(img[111]), .B1(n28433), .B2(n30197), .O(
        n24453) );
  ND2S U25983 ( .I1(n24340), .I2(n24453), .O(n24454) );
  NR2 U25984 ( .I1(n24023), .I2(n24957), .O(n29027) );
  AOI22S U25985 ( .A1(n13772), .A2(img[1239]), .B1(n28862), .B2(n30198), .O(
        n24455) );
  ND2S U25986 ( .I1(n24340), .I2(n24455), .O(n24456) );
  AOI22S U25987 ( .A1(n28614), .A2(n30199), .B1(n24808), .B2(img[1199]), .O(
        n24458) );
  ND3S U25988 ( .I1(n24340), .I2(n24458), .I3(n24457), .O(n24459) );
  MUX2 U25989 ( .A(img[1239]), .B(n24459), .S(n29037), .O(n12293) );
  AOI22S U25990 ( .A1(n28162), .A2(n30200), .B1(n24808), .B2(img[1175]), .O(
        n24461) );
  ND3S U25991 ( .I1(n24340), .I2(n24461), .I3(n24460), .O(n24464) );
  MUX2 U25992 ( .A(img[1263]), .B(n24464), .S(n29044), .O(n12275) );
  AOI22S U25993 ( .A1(n28347), .A2(img[1263]), .B1(n23941), .B2(n30201), .O(
        n24465) );
  ND2S U25994 ( .I1(n24340), .I2(n24465), .O(n24467) );
  AOI22S U25995 ( .A1(n26101), .A2(img[1367]), .B1(n23918), .B2(n30202), .O(
        n24468) );
  ND2S U25996 ( .I1(n24340), .I2(n24468), .O(n24470) );
  MUX2 U25997 ( .A(n24470), .B(img[1327]), .S(n29047), .O(n12205) );
  AOI22S U25998 ( .A1(n29096), .A2(n30203), .B1(n24808), .B2(img[1327]), .O(
        n24472) );
  ND3S U25999 ( .I1(n24340), .I2(n24472), .I3(n24471), .O(n24473) );
  MUX2 U26000 ( .A(img[1367]), .B(n24473), .S(n29051), .O(n12171) );
  AOI22S U26001 ( .A1(n29096), .A2(n30204), .B1(n24808), .B2(img[1303]), .O(
        n24475) );
  ND3S U26002 ( .I1(n24340), .I2(n24475), .I3(n24474), .O(n24477) );
  MUX2 U26003 ( .A(img[1391]), .B(n24477), .S(n29058), .O(n12141) );
  AOI22S U26004 ( .A1(n13771), .A2(img[1391]), .B1(n13779), .B2(n30205), .O(
        n24478) );
  ND2S U26005 ( .I1(n24340), .I2(n24478), .O(n24480) );
  MUX2 U26006 ( .A(n24480), .B(img[1303]), .S(n29054), .O(n12235) );
  AOI22S U26007 ( .A1(n25810), .A2(img[919]), .B1(n27511), .B2(n30206), .O(
        n24481) );
  ND2S U26008 ( .I1(n24340), .I2(n24481), .O(n24483) );
  NR2 U26009 ( .I1(n24542), .I2(n24716), .O(n24482) );
  NR2P U26010 ( .I1(n24482), .I2(n24717), .O(n29064) );
  AOI22S U26011 ( .A1(n28106), .A2(img[1007]), .B1(n24193), .B2(n30207), .O(
        n24484) );
  ND2S U26012 ( .I1(n24340), .I2(n24484), .O(n24485) );
  OAI12HS U26013 ( .B1(n24023), .B2(n24713), .A1(n24495), .O(n29061) );
  MUX2 U26014 ( .A(img[919]), .B(n24485), .S(n29061), .O(n12613) );
  AOI22S U26015 ( .A1(n28347), .A2(img[151]), .B1(n28913), .B2(n30208), .O(
        n24486) );
  ND2S U26016 ( .I1(n24340), .I2(n24486), .O(n24488) );
  INV1S U26017 ( .I(n24529), .O(n24487) );
  MUX2 U26018 ( .A(img[239]), .B(n24488), .S(n29070), .O(n13299) );
  AOI22S U26019 ( .A1(n26970), .A2(img[239]), .B1(n29407), .B2(n30209), .O(
        n24489) );
  ND2S U26020 ( .I1(n24340), .I2(n24489), .O(n24491) );
  MUX2 U26021 ( .A(img[151]), .B(n24491), .S(n29067), .O(n13381) );
  AOI22S U26022 ( .A1(n13772), .A2(img[279]), .B1(n28695), .B2(n30210), .O(
        n24492) );
  ND2S U26023 ( .I1(n24340), .I2(n24492), .O(n24493) );
  OAI12HS U26024 ( .B1(n24732), .B2(n24529), .A1(n24495), .O(n29078) );
  MUX2 U26025 ( .A(img[367]), .B(n24493), .S(n29078), .O(n13165) );
  AOI22S U26026 ( .A1(n13780), .A2(img[367]), .B1(n24755), .B2(n30211), .O(
        n24494) );
  ND2S U26027 ( .I1(n24340), .I2(n24494), .O(n24496) );
  OAI12HS U26028 ( .B1(n24732), .B2(n24023), .A1(n24495), .O(n29074) );
  AOI22S U26029 ( .A1(n29414), .A2(img[407]), .B1(n25591), .B2(n30212), .O(
        n24497) );
  ND2S U26030 ( .I1(n24340), .I2(n24497), .O(n24498) );
  MUX2 U26031 ( .A(img[495]), .B(n24498), .S(n29084), .O(n13043) );
  AOI22S U26032 ( .A1(n28347), .A2(img[495]), .B1(n25377), .B2(n30213), .O(
        n24499) );
  ND2S U26033 ( .I1(n24340), .I2(n24499), .O(n24502) );
  AOI22S U26034 ( .A1(n29435), .A2(img[1495]), .B1(n27735), .B2(n30214), .O(
        n24503) );
  ND2S U26035 ( .I1(n24340), .I2(n24503), .O(n24505) );
  ND2S U26036 ( .I1(n24758), .I2(n24520), .O(n24504) );
  ND2 U26037 ( .I1(n24590), .I2(n24504), .O(n29087) );
  MUX2 U26038 ( .A(n24505), .B(img[1455]), .S(n29087), .O(n12083) );
  AOI22S U26039 ( .A1(n13779), .A2(n30215), .B1(n24808), .B2(img[1455]), .O(
        n24507) );
  INV1S U26040 ( .I(n24585), .O(n24508) );
  NR2 U26041 ( .I1(n24509), .I2(n24508), .O(n24511) );
  AOI22S U26042 ( .A1(n13779), .A2(n30216), .B1(n24808), .B2(img[1431]), .O(
        n24514) );
  ND3S U26043 ( .I1(n24340), .I2(n24514), .I3(n24513), .O(n24518) );
  MUX2 U26044 ( .A(img[1519]), .B(n24518), .S(n29099), .O(n12019) );
  AOI22S U26045 ( .A1(n27722), .A2(img[1519]), .B1(n27735), .B2(n30217), .O(
        n24519) );
  ND2S U26046 ( .I1(n24340), .I2(n24519), .O(n24521) );
  OAI12HS U26047 ( .B1(n24023), .B2(n24520), .A1(n24495), .O(n29094) );
  INV1S U26048 ( .I(img[879]), .O(n24522) );
  AOI22S U26049 ( .A1(n25810), .A2(img[791]), .B1(n13775), .B2(n24522), .O(
        n24523) );
  ND2S U26050 ( .I1(n24340), .I2(n24523), .O(n24525) );
  ND2S U26051 ( .I1(n24748), .I2(n24529), .O(n24524) );
  AOI22S U26052 ( .A1(n27722), .A2(img[879]), .B1(n28862), .B2(n30218), .O(
        n24526) );
  ND2S U26053 ( .I1(n24340), .I2(n24526), .O(n24527) );
  OAI12HS U26054 ( .B1(n24023), .B2(n24744), .A1(n24495), .O(n29102) );
  MUX2 U26055 ( .A(img[791]), .B(n24527), .S(n29102), .O(n12747) );
  AOI22S U26056 ( .A1(n27722), .A2(img[663]), .B1(n27049), .B2(n30219), .O(
        n24528) );
  ND2S U26057 ( .I1(n24424), .I2(n24528), .O(n24531) );
  ND2S U26058 ( .I1(n24758), .I2(n24529), .O(n24530) );
  MUX2 U26059 ( .A(n24531), .B(img[751]), .S(n29112), .O(n12787) );
  AOI22S U26060 ( .A1(n13773), .A2(img[751]), .B1(n29457), .B2(n30220), .O(
        n24532) );
  ND2S U26061 ( .I1(n24340), .I2(n24532), .O(n24533) );
  OAI12HS U26062 ( .B1(n24023), .B2(n24753), .A1(n24495), .O(n29109) );
  AOI22S U26063 ( .A1(n27110), .A2(img[1111]), .B1(n29397), .B2(n30221), .O(
        n24534) );
  ND2S U26064 ( .I1(n24340), .I2(n24534), .O(n24535) );
  MUX2 U26065 ( .A(n24535), .B(img[1071]), .S(n29115), .O(n12461) );
  AOI22S U26066 ( .A1(n28037), .A2(n30222), .B1(n24808), .B2(img[1071]), .O(
        n24537) );
  ND2S U26067 ( .I1(n13770), .I2(img[1135]), .O(n24536) );
  ND3S U26068 ( .I1(n24340), .I2(n24537), .I3(n24536), .O(n24538) );
  MUX2 U26069 ( .A(img[1111]), .B(n24538), .S(n29119), .O(n12427) );
  AOI22S U26070 ( .A1(n28343), .A2(n30223), .B1(n24808), .B2(img[1047]), .O(
        n24540) );
  ND3S U26071 ( .I1(n24340), .I2(n24540), .I3(n24539), .O(n24544) );
  MUX2 U26072 ( .A(img[1135]), .B(n24544), .S(n29127), .O(n12397) );
  AOI22S U26073 ( .A1(n29072), .A2(img[1135]), .B1(n28913), .B2(n30224), .O(
        n24545) );
  ND2S U26074 ( .I1(n24340), .I2(n24545), .O(n24547) );
  MUX2 U26075 ( .A(n24547), .B(img[1047]), .S(n29122), .O(n12490) );
  AOI22S U26076 ( .A1(n13773), .A2(img[559]), .B1(n29407), .B2(n30225), .O(
        n24548) );
  ND2S U26077 ( .I1(n24340), .I2(n24548), .O(n24549) );
  NR2 U26078 ( .I1(n24585), .I2(n24692), .O(n24578) );
  AO12 U26079 ( .B1(n24578), .B2(n24694), .A1(n24693), .O(n29133) );
  MUX2 U26080 ( .A(n24549), .B(img[599]), .S(n29133), .O(n12939) );
  AOI22S U26081 ( .A1(n26970), .A2(img[599]), .B1(n29457), .B2(n30226), .O(
        n24550) );
  ND2S U26082 ( .I1(n24340), .I2(n24550), .O(n24551) );
  AO12 U26083 ( .B1(n24563), .B2(n24694), .A1(n24693), .O(n29439) );
  MUX2 U26084 ( .A(n24551), .B(img[559]), .S(n29439), .O(n12973) );
  AOI22S U26085 ( .A1(n28442), .A2(img[47]), .B1(n25591), .B2(n30227), .O(
        n24552) );
  ND2S U26086 ( .I1(n24340), .I2(n24552), .O(n24553) );
  AOI22S U26087 ( .A1(n26490), .A2(img[87]), .B1(n29397), .B2(n30228), .O(
        n24554) );
  ND2S U26088 ( .I1(n24340), .I2(n24554), .O(n24555) );
  MUX2 U26089 ( .A(img[47]), .B(n24555), .S(n29136), .O(n13485) );
  AOI22S U26090 ( .A1(n27685), .A2(img[175]), .B1(n25591), .B2(n30229), .O(
        n24556) );
  ND2S U26091 ( .I1(n24340), .I2(n24556), .O(n24557) );
  MUX2 U26092 ( .A(img[215]), .B(n24557), .S(n29151), .O(n13317) );
  AOI22S U26093 ( .A1(n28347), .A2(img[215]), .B1(n28913), .B2(n30230), .O(
        n24558) );
  ND2S U26094 ( .I1(n24340), .I2(n24558), .O(n24559) );
  MUX2 U26095 ( .A(img[175]), .B(n24559), .S(n29148), .O(n13363) );
  AOI22S U26096 ( .A1(n25595), .A2(img[303]), .B1(n28938), .B2(n30231), .O(
        n24560) );
  ND2S U26097 ( .I1(n24340), .I2(n24560), .O(n24561) );
  OAI12HS U26098 ( .B1(n24732), .B2(n24578), .A1(n24495), .O(n29157) );
  AOI22S U26099 ( .A1(n26101), .A2(img[343]), .B1(n28695), .B2(n30232), .O(
        n24562) );
  ND2S U26100 ( .I1(n24340), .I2(n24562), .O(n24564) );
  OAI12HS U26101 ( .B1(n24732), .B2(n24563), .A1(n24495), .O(n29154) );
  MUX2 U26102 ( .A(img[303]), .B(n24564), .S(n29154), .O(n13229) );
  AOI22S U26103 ( .A1(n27722), .A2(img[431]), .B1(n24374), .B2(n30233), .O(
        n24565) );
  ND2S U26104 ( .I1(n24340), .I2(n24565), .O(n24566) );
  MUX2 U26105 ( .A(img[471]), .B(n24566), .S(n29163), .O(n13061) );
  AOI22S U26106 ( .A1(n27722), .A2(img[471]), .B1(n29194), .B2(n30234), .O(
        n24567) );
  ND2S U26107 ( .I1(n24340), .I2(n24567), .O(n24569) );
  OA12 U26108 ( .B1(n24568), .B2(n24669), .A1(n24668), .O(n29160) );
  MUX2 U26109 ( .A(img[431]), .B(n24569), .S(n29160), .O(n13107) );
  INV1S U26110 ( .I(img[855]), .O(n24570) );
  AOI22S U26111 ( .A1(n13773), .A2(img[815]), .B1(n28075), .B2(n24570), .O(
        n24571) );
  ND2S U26112 ( .I1(n24340), .I2(n24571), .O(n24573) );
  ND2S U26113 ( .I1(n24748), .I2(n24578), .O(n24572) );
  AOI22S U26114 ( .A1(n27722), .A2(img[855]), .B1(n28862), .B2(n30235), .O(
        n24574) );
  ND2S U26115 ( .I1(n24340), .I2(n24574), .O(n24576) );
  MUX2 U26116 ( .A(n24576), .B(img[815]), .S(n29166), .O(n12717) );
  AOI22S U26117 ( .A1(n26822), .A2(img[687]), .B1(n24374), .B2(n30236), .O(
        n24577) );
  ND2S U26118 ( .I1(n24340), .I2(n24577), .O(n24580) );
  ND2S U26119 ( .I1(n24758), .I2(n24578), .O(n24579) );
  BUF2 U26120 ( .I(n24581), .O(n24658) );
  AOI22S U26121 ( .A1(n27722), .A2(img[727]), .B1(n24374), .B2(n30237), .O(
        n24582) );
  ND2S U26122 ( .I1(n24658), .I2(n24582), .O(n24583) );
  AOI22S U26123 ( .A1(n27722), .A2(img[943]), .B1(n28075), .B2(n30238), .O(
        n24584) );
  ND2S U26124 ( .I1(n24658), .I2(n24584), .O(n24587) );
  NR2 U26125 ( .I1(n24585), .I2(n24716), .O(n24586) );
  NR2P U26126 ( .I1(n24586), .I2(n24717), .O(n29145) );
  MUX2 U26127 ( .A(img[983]), .B(n24587), .S(n29145), .O(n12549) );
  AOI22S U26128 ( .A1(n27746), .A2(img[983]), .B1(n28075), .B2(n30239), .O(
        n24588) );
  ND2S U26129 ( .I1(n24658), .I2(n24588), .O(n24591) );
  ND2S U26130 ( .I1(n24758), .I2(n24713), .O(n24589) );
  AOI22S U26131 ( .A1(n27746), .A2(img[351]), .B1(n25062), .B2(n30240), .O(
        n24592) );
  ND2S U26132 ( .I1(n24658), .I2(n24592), .O(n24593) );
  OAI12HS U26133 ( .B1(n24732), .B2(n24612), .A1(n24495), .O(n29361) );
  AOI22S U26134 ( .A1(n27746), .A2(img[295]), .B1(n28433), .B2(n30241), .O(
        n24594) );
  ND2S U26135 ( .I1(n24658), .I2(n24594), .O(n24595) );
  NR2 U26136 ( .I1(n24622), .I2(n24692), .O(n24636) );
  OAI12HS U26137 ( .B1(n24732), .B2(n24636), .A1(n24495), .O(n29358) );
  MUX2 U26138 ( .A(img[351]), .B(n24595), .S(n29358), .O(n13181) );
  AOI22S U26139 ( .A1(n27746), .A2(img[607]), .B1(n13781), .B2(n30242), .O(
        n24596) );
  ND2S U26140 ( .I1(n24658), .I2(n24596), .O(n24598) );
  INV1S U26141 ( .I(n24693), .O(n24597) );
  AOI22S U26142 ( .A1(n28347), .A2(img[551]), .B1(n25591), .B2(n30243), .O(
        n24599) );
  ND2S U26143 ( .I1(n24658), .I2(n24599), .O(n24600) );
  AO12 U26144 ( .B1(n24636), .B2(n24694), .A1(n24693), .O(n29478) );
  MUX2 U26145 ( .A(n24600), .B(img[607]), .S(n29478), .O(n12925) );
  AOI22S U26146 ( .A1(n29414), .A2(img[95]), .B1(n28037), .B2(n30244), .O(
        n24601) );
  ND2S U26147 ( .I1(n24658), .I2(n24601), .O(n24602) );
  MUX2 U26148 ( .A(img[39]), .B(n24602), .S(n29342), .O(n13499) );
  AOI22S U26149 ( .A1(n28382), .A2(img[39]), .B1(n29530), .B2(n30245), .O(
        n24603) );
  ND2S U26150 ( .I1(n24658), .I2(n24603), .O(n24604) );
  MUX2 U26151 ( .A(img[95]), .B(n24604), .S(n29339), .O(n13437) );
  AOI22S U26152 ( .A1(n29129), .A2(img[991]), .B1(n23941), .B2(n30246), .O(
        n24605) );
  ND2S U26153 ( .I1(n24658), .I2(n24605), .O(n24607) );
  ND2S U26154 ( .I1(n24713), .I2(n24694), .O(n24606) );
  AOI22S U26155 ( .A1(n27685), .A2(img[935]), .B1(n27049), .B2(n30247), .O(
        n24608) );
  ND2S U26156 ( .I1(n24658), .I2(n24608), .O(n24610) );
  NR2 U26157 ( .I1(n24622), .I2(n24716), .O(n24609) );
  NR2P U26158 ( .I1(n24609), .I2(n24717), .O(n29345) );
  MUX2 U26159 ( .A(img[991]), .B(n24610), .S(n29345), .O(n12547) );
  AOI22S U26160 ( .A1(n27685), .A2(img[223]), .B1(n13781), .B2(n30248), .O(
        n24611) );
  ND2S U26161 ( .I1(n24658), .I2(n24611), .O(n24615) );
  INV1S U26162 ( .I(n24612), .O(n24613) );
  MUX2 U26163 ( .A(img[167]), .B(n24615), .S(n29355), .O(n13365) );
  AOI22S U26164 ( .A1(n25810), .A2(img[167]), .B1(n25377), .B2(n30249), .O(
        n24616) );
  ND2S U26165 ( .I1(n24658), .I2(n24616), .O(n24617) );
  MUX2 U26166 ( .A(img[223]), .B(n24617), .S(n29351), .O(n13315) );
  AOI22S U26167 ( .A1(n25595), .A2(img[479]), .B1(n27049), .B2(n30250), .O(
        n24618) );
  ND2S U26168 ( .I1(n24658), .I2(n24618), .O(n24620) );
  OA12 U26169 ( .B1(n24619), .B2(n24669), .A1(n24668), .O(n29367) );
  MUX2 U26170 ( .A(img[423]), .B(n24620), .S(n29367), .O(n13109) );
  AOI22S U26171 ( .A1(n25595), .A2(img[423]), .B1(n25591), .B2(n30251), .O(
        n24621) );
  ND2S U26172 ( .I1(n24658), .I2(n24621), .O(n24623) );
  MUX2 U26173 ( .A(img[479]), .B(n24623), .S(n29364), .O(n13059) );
  AOI22S U26174 ( .A1(n28083), .A2(img[863]), .B1(n25591), .B2(n30252), .O(
        n24624) );
  ND2S U26175 ( .I1(n24658), .I2(n24624), .O(n24626) );
  MUX2 U26176 ( .A(n24626), .B(img[807]), .S(n29374), .O(n12731) );
  INV1S U26177 ( .I(img[863]), .O(n24627) );
  AOI22S U26178 ( .A1(n25810), .A2(img[807]), .B1(n28695), .B2(n24627), .O(
        n24628) );
  ND2S U26179 ( .I1(n24658), .I2(n24628), .O(n24630) );
  ND2S U26180 ( .I1(n24748), .I2(n24636), .O(n24629) );
  AOI22S U26181 ( .A1(n27746), .A2(img[735]), .B1(n13781), .B2(n30253), .O(
        n24631) );
  ND2S U26182 ( .I1(n24658), .I2(n24631), .O(n24634) );
  ND2S U26183 ( .I1(n24753), .I2(n24694), .O(n24632) );
  AOI22S U26184 ( .A1(n27746), .A2(img[679]), .B1(n13781), .B2(n30254), .O(
        n24635) );
  ND2S U26185 ( .I1(n24658), .I2(n24635), .O(n24638) );
  ND2S U26186 ( .I1(n24758), .I2(n24636), .O(n24637) );
  MUX2 U26187 ( .A(n24638), .B(img[735]), .S(n29377), .O(n12803) );
  AOI22S U26188 ( .A1(n27746), .A2(img[631]), .B1(n24374), .B2(n30255), .O(
        n24639) );
  ND2S U26189 ( .I1(n24658), .I2(n24639), .O(n24642) );
  NR2 U26190 ( .I1(n24640), .I2(n24726), .O(n24641) );
  AOI22S U26191 ( .A1(n27746), .A2(img[527]), .B1(n24374), .B2(n30256), .O(
        n24643) );
  ND2S U26192 ( .I1(n24658), .I2(n24643), .O(n24644) );
  NR2 U26193 ( .I1(n24670), .I2(n24692), .O(n24958) );
  AO12 U26194 ( .B1(n24958), .B2(n24694), .A1(n24693), .O(n29292) );
  MUX2 U26195 ( .A(n24644), .B(img[631]), .S(n29292), .O(n12907) );
  AOI22S U26196 ( .A1(n27746), .A2(img[1015]), .B1(n29457), .B2(n30257), .O(
        n24645) );
  ND2S U26197 ( .I1(n24658), .I2(n24645), .O(n24648) );
  NR2 U26198 ( .I1(n24646), .I2(n24726), .O(n24647) );
  AOI22S U26199 ( .A1(n27746), .A2(img[911]), .B1(n28862), .B2(n30258), .O(
        n24649) );
  ND2S U26200 ( .I1(n24658), .I2(n24649), .O(n24651) );
  NR2 U26201 ( .I1(n24670), .I2(n24716), .O(n24650) );
  NR2P U26202 ( .I1(n24650), .I2(n24717), .O(n29303) );
  MUX2 U26203 ( .A(img[1015]), .B(n24651), .S(n29303), .O(n12517) );
  AOI22S U26204 ( .A1(n27746), .A2(img[247]), .B1(n25591), .B2(n30259), .O(
        n24652) );
  ND2S U26205 ( .I1(n24658), .I2(n24652), .O(n24654) );
  INV1S U26206 ( .I(n24725), .O(n24653) );
  AOI22S U26207 ( .A1(n27990), .A2(img[143]), .B1(n24374), .B2(n30260), .O(
        n24655) );
  ND2S U26208 ( .I1(n24658), .I2(n24655), .O(n24656) );
  MUX2 U26209 ( .A(img[247]), .B(n24656), .S(n29309), .O(n13285) );
  AOI22S U26210 ( .A1(n28347), .A2(img[375]), .B1(n28862), .B2(n30261), .O(
        n24657) );
  ND2S U26211 ( .I1(n24658), .I2(n24657), .O(n24660) );
  MUX2 U26212 ( .A(n24660), .B(img[271]), .S(n29312), .O(n13261) );
  AOI22S U26213 ( .A1(n25810), .A2(img[271]), .B1(n28913), .B2(n30262), .O(
        n24661) );
  ND2S U26214 ( .I1(n24340), .I2(n24661), .O(n24662) );
  OAI12HS U26215 ( .B1(n24732), .B2(n24958), .A1(n24495), .O(n29315) );
  AOI22S U26216 ( .A1(n28442), .A2(img[503]), .B1(n13781), .B2(n30263), .O(
        n24663) );
  ND2S U26217 ( .I1(n24340), .I2(n24663), .O(n24666) );
  AOI22S U26218 ( .A1(n24415), .A2(img[399]), .B1(n25062), .B2(n30264), .O(
        n24667) );
  ND2S U26219 ( .I1(n24340), .I2(n24667), .O(n24671) );
  MUX2 U26220 ( .A(img[503]), .B(n24671), .S(n29321), .O(n13029) );
  AOI22S U26221 ( .A1(n27065), .A2(img[887]), .B1(n29194), .B2(n30265), .O(
        n24672) );
  ND2S U26222 ( .I1(n24340), .I2(n24672), .O(n24675) );
  NR2 U26223 ( .I1(n24673), .I2(n24726), .O(n24674) );
  MUX2 U26224 ( .A(img[783]), .B(n24675), .S(n29324), .O(n12749) );
  INV1S U26225 ( .I(img[887]), .O(n24676) );
  AOI22S U26226 ( .A1(n13778), .A2(img[783]), .B1(n28135), .B2(n24676), .O(
        n24677) );
  ND2S U26227 ( .I1(n24340), .I2(n24677), .O(n24679) );
  ND2S U26228 ( .I1(n24748), .I2(n24958), .O(n24678) );
  AOI22S U26229 ( .A1(n28318), .A2(img[759]), .B1(n25062), .B2(n30266), .O(
        n24680) );
  ND2S U26230 ( .I1(n24340), .I2(n24680), .O(n24684) );
  NR2 U26231 ( .I1(n24681), .I2(n24726), .O(n24683) );
  AOI22S U26232 ( .A1(n27110), .A2(img[655]), .B1(n28614), .B2(n30267), .O(
        n24685) );
  ND2S U26233 ( .I1(n24340), .I2(n24685), .O(n24687) );
  ND2S U26234 ( .I1(n24758), .I2(n24958), .O(n24686) );
  AOI22S U26235 ( .A1(n27065), .A2(img[639]), .B1(n28862), .B2(n30268), .O(
        n24688) );
  ND2S U26236 ( .I1(n24340), .I2(n24688), .O(n24690) );
  INV1S U26237 ( .I(n24229), .O(n24736) );
  AOI22S U26238 ( .A1(n29414), .A2(img[519]), .B1(n28433), .B2(n30269), .O(
        n24691) );
  ND2S U26239 ( .I1(n24340), .I2(n24691), .O(n24695) );
  NR2 U26240 ( .I1(n24727), .I2(n24692), .O(n24757) );
  AO12 U26241 ( .B1(n24757), .B2(n24694), .A1(n24693), .O(n29386) );
  MUX2 U26242 ( .A(n24695), .B(img[639]), .S(n29386), .O(n12893) );
  AOI22S U26243 ( .A1(n28468), .A2(img[127]), .B1(n25062), .B2(n30270), .O(
        n24696) );
  ND2S U26244 ( .I1(n24340), .I2(n24696), .O(n24709) );
  INV1S U26245 ( .I(n24697), .O(n24765) );
  OAI22S U26246 ( .A1(n24701), .A2(n24700), .B1(n24699), .B2(n24698), .O(
        n24704) );
  NR3 U26247 ( .I1(n24706), .I2(n24702), .I3(n28575), .O(n24703) );
  NR2 U26248 ( .I1(n24704), .I2(n24703), .O(n24707) );
  AOI13HS U26249 ( .B1(n24765), .B2(n24708), .B3(n24764), .A1(n24763), .O(
        n29389) );
  AOI22S U26250 ( .A1(n28468), .A2(img[7]), .B1(n13781), .B2(n30271), .O(
        n24710) );
  ND2S U26251 ( .I1(n24340), .I2(n24710), .O(n24711) );
  MUX2 U26252 ( .A(img[127]), .B(n24711), .S(n29392), .O(n13405) );
  AOI22S U26253 ( .A1(n28468), .A2(img[1023]), .B1(n28075), .B2(n30272), .O(
        n24712) );
  ND2S U26254 ( .I1(n24340), .I2(n24712), .O(n24714) );
  MUX2 U26255 ( .A(img[903]), .B(n24714), .S(n29395), .O(n12629) );
  AOI22S U26256 ( .A1(n28468), .A2(img[903]), .B1(n13781), .B2(n30273), .O(
        n24715) );
  ND2S U26257 ( .I1(n24340), .I2(n24715), .O(n24719) );
  NR2 U26258 ( .I1(n24727), .I2(n24716), .O(n24718) );
  NR2P U26259 ( .I1(n24718), .I2(n24717), .O(n29399) );
  AOI22S U26260 ( .A1(n27722), .A2(img[255]), .B1(n28913), .B2(n30274), .O(
        n24720) );
  ND2S U26261 ( .I1(n24340), .I2(n24720), .O(n24723) );
  MUX2 U26262 ( .A(n24723), .B(img[135]), .S(n29402), .O(n13397) );
  AOI22S U26263 ( .A1(n26101), .A2(img[135]), .B1(n24193), .B2(n30275), .O(
        n24724) );
  ND2S U26264 ( .I1(n24340), .I2(n24724), .O(n24728) );
  MUX2 U26265 ( .A(img[255]), .B(n24728), .S(n29405), .O(n13282) );
  AOI22S U26266 ( .A1(n26101), .A2(img[383]), .B1(n23941), .B2(n30276), .O(
        n24729) );
  ND2S U26267 ( .I1(n24340), .I2(n24729), .O(n24730) );
  AOI22S U26268 ( .A1(n25595), .A2(img[263]), .B1(n13781), .B2(n30277), .O(
        n24731) );
  ND2S U26269 ( .I1(n24340), .I2(n24731), .O(n24733) );
  OAI12HS U26270 ( .B1(n24732), .B2(n24757), .A1(n24495), .O(n29412) );
  MUX2 U26271 ( .A(img[383]), .B(n24733), .S(n29412), .O(n13149) );
  AOI22S U26272 ( .A1(n28347), .A2(img[511]), .B1(n28162), .B2(n30278), .O(
        n24734) );
  ND2S U26273 ( .I1(n24340), .I2(n24734), .O(n24737) );
  MUX2 U26274 ( .A(n24737), .B(img[391]), .S(n29416), .O(n13141) );
  INV1S U26275 ( .I(img[511]), .O(n24738) );
  AOI22S U26276 ( .A1(n25810), .A2(img[391]), .B1(n28938), .B2(n24738), .O(
        n24739) );
  ND2S U26277 ( .I1(n24340), .I2(n24739), .O(n24742) );
  AO12 U26278 ( .B1(n24757), .B2(n24741), .A1(n24740), .O(n29420) );
  AOI22S U26279 ( .A1(n27957), .A2(img[895]), .B1(n25062), .B2(n30279), .O(
        n24743) );
  ND2S U26280 ( .I1(n24340), .I2(n24743), .O(n24745) );
  MUX2 U26281 ( .A(img[775]), .B(n24745), .S(n29423), .O(n12763) );
  INV1S U26282 ( .I(img[895]), .O(n24746) );
  AOI22S U26283 ( .A1(n28347), .A2(img[775]), .B1(n13781), .B2(n24746), .O(
        n24747) );
  ND2S U26284 ( .I1(n24340), .I2(n24747), .O(n24751) );
  ND2S U26285 ( .I1(n24748), .I2(n24757), .O(n24749) );
  AOI22S U26286 ( .A1(n29072), .A2(img[767]), .B1(n29194), .B2(n30280), .O(
        n24752) );
  ND2S U26287 ( .I1(n24340), .I2(n24752), .O(n24754) );
  AOI22S U26288 ( .A1(n27065), .A2(img[647]), .B1(n25859), .B2(n30281), .O(
        n24756) );
  ND2S U26289 ( .I1(n24340), .I2(n24756), .O(n24761) );
  ND2S U26290 ( .I1(n24758), .I2(n24757), .O(n24759) );
  AOI22S U26291 ( .A1(n26970), .A2(img[119]), .B1(n28862), .B2(n30282), .O(
        n24762) );
  ND2S U26292 ( .I1(n24340), .I2(n24762), .O(n24767) );
  AOI13HS U26293 ( .B1(n24766), .B2(n24765), .B3(n24764), .A1(n24763), .O(
        n29295) );
  INV1S U26294 ( .I(n21416), .O(n24772) );
  OAI22S U26295 ( .A1(n24769), .A2(n28530), .B1(n13897), .B2(n24768), .O(
        n24770) );
  OAI12HS U26296 ( .B1(n28536), .B2(n24772), .A1(n24771), .O(n24794) );
  INV1S U26297 ( .I(A67_shift[46]), .O(n24775) );
  AOI22S U26298 ( .A1(n28553), .A2(A67_shift[14]), .B1(n28546), .B2(
        A67_shift[174]), .O(n24774) );
  AOI12HS U26299 ( .B1(n28552), .B2(A67_shift[142]), .A1(n28540), .O(n24773)
         );
  OAI112HS U26300 ( .C1(n28544), .C2(n24775), .A1(n24774), .B1(n24773), .O(
        n24788) );
  ND2S U26301 ( .I1(n28547), .I2(A67_shift[238]), .O(n24778) );
  AOI22S U26302 ( .A1(n28550), .A2(A67_shift[78]), .B1(n28551), .B2(
        A67_shift[206]), .O(n24777) );
  ND2S U26303 ( .I1(n28554), .I2(A67_shift[110]), .O(n24776) );
  ND2S U26304 ( .I1(n28547), .I2(A67_shift[254]), .O(n24781) );
  AOI22S U26305 ( .A1(n28552), .A2(A67_shift[158]), .B1(n28551), .B2(
        A67_shift[222]), .O(n24780) );
  ND2S U26306 ( .I1(n28554), .I2(A67_shift[126]), .O(n24779) );
  INV1S U26307 ( .I(A67_shift[62]), .O(n24784) );
  AOI22S U26308 ( .A1(n28553), .A2(A67_shift[30]), .B1(n28546), .B2(
        A67_shift[190]), .O(n24783) );
  AOI12HS U26309 ( .B1(n28550), .B2(A67_shift[94]), .A1(n28555), .O(n24782) );
  OAI112HS U26310 ( .C1(n28544), .C2(n24784), .A1(n24783), .B1(n24782), .O(
        n24785) );
  OAI22S U26311 ( .A1(n24788), .A2(n24787), .B1(n24786), .B2(n24785), .O(
        n24792) );
  AOI22S U26312 ( .A1(n28566), .A2(gray_max_out[6]), .B1(n28565), .B2(
        gray_weight_out[6]), .O(n24790) );
  ND2S U26313 ( .I1(n28564), .I2(gray_avg_out[6]), .O(n24789) );
  AOI12HT U26314 ( .B1(n24794), .B2(n28575), .A1(n24793), .O(n25298) );
  AOI22S U26315 ( .A1(n26101), .A2(img[574]), .B1(n28135), .B2(n30283), .O(
        n24795) );
  ND2S U26316 ( .I1(n25327), .I2(n24795), .O(n24796) );
  MUX2 U26317 ( .A(n24796), .B(img[582]), .S(n28799), .O(n12954) );
  AOI22S U26318 ( .A1(n28468), .A2(img[70]), .B1(n25591), .B2(n30284), .O(
        n24797) );
  ND2S U26319 ( .I1(n25327), .I2(n24797), .O(n24798) );
  AOI22S U26320 ( .A1(n28468), .A2(img[62]), .B1(n28695), .B2(n30285), .O(
        n24799) );
  ND2S U26321 ( .I1(n25327), .I2(n24799), .O(n24800) );
  MUX2 U26322 ( .A(img[70]), .B(n24800), .S(n28804), .O(n13466) );
  AOI22S U26323 ( .A1(n28468), .A2(img[1278]), .B1(n13781), .B2(n30286), .O(
        n24801) );
  ND2S U26324 ( .I1(n25327), .I2(n24801), .O(n24802) );
  AOI22S U26325 ( .A1(n28913), .A2(n30287), .B1(n24808), .B2(img[1158]), .O(
        n24804) );
  ND2S U26326 ( .I1(n13770), .I2(img[1222]), .O(n24803) );
  ND3S U26327 ( .I1(n25327), .I2(n24804), .I3(n24803), .O(n24805) );
  MUX2 U26328 ( .A(img[1278]), .B(n24805), .S(n28814), .O(n12258) );
  AOI22S U26329 ( .A1(n28468), .A2(img[1222]), .B1(n28592), .B2(n30288), .O(
        n24806) );
  ND2S U26330 ( .I1(n25327), .I2(n24806), .O(n24807) );
  MUX2 U26331 ( .A(img[1214]), .B(n24807), .S(n28821), .O(n12322) );
  AOI22S U26332 ( .A1(n27049), .A2(n30289), .B1(n24808), .B2(img[1214]), .O(
        n24810) );
  ND2S U26333 ( .I1(n13902), .I2(img[1278]), .O(n24809) );
  ND3S U26334 ( .I1(n25327), .I2(n24810), .I3(n24809), .O(n24811) );
  MUX2 U26335 ( .A(img[1222]), .B(n24811), .S(n28818), .O(n12310) );
  AOI22S U26336 ( .A1(n28468), .A2(img[1406]), .B1(n29242), .B2(n30290), .O(
        n24812) );
  ND2S U26337 ( .I1(n25327), .I2(n24812), .O(n24813) );
  MUX2 U26338 ( .A(img[1286]), .B(n24813), .S(n28824), .O(n12250) );
  AOI22S U26339 ( .A1(n25468), .A2(n30291), .B1(n24890), .B2(img[1286]), .O(
        n24815) );
  ND3S U26340 ( .I1(n25327), .I2(n24815), .I3(n24814), .O(n24816) );
  MUX2 U26341 ( .A(img[1406]), .B(n24816), .S(n28828), .O(n12126) );
  AOI22S U26342 ( .A1(n28468), .A2(img[1350]), .B1(n27049), .B2(n30292), .O(
        n24817) );
  ND2S U26343 ( .I1(n25327), .I2(n24817), .O(n24818) );
  AOI22S U26344 ( .A1(n25377), .A2(n30293), .B1(n24890), .B2(img[1342]), .O(
        n24820) );
  ND3S U26345 ( .I1(n25327), .I2(n24820), .I3(n24819), .O(n24821) );
  MUX2 U26346 ( .A(img[1350]), .B(n24821), .S(n28832), .O(n12186) );
  AOI22S U26347 ( .A1(n28083), .A2(img[966]), .B1(n25591), .B2(n30294), .O(
        n24822) );
  ND2S U26348 ( .I1(n25327), .I2(n24822), .O(n24823) );
  MUX2 U26349 ( .A(img[958]), .B(n24823), .S(n28842), .O(n12578) );
  AOI22S U26350 ( .A1(n27746), .A2(img[958]), .B1(n25062), .B2(n30295), .O(
        n24824) );
  ND2S U26351 ( .I1(n25327), .I2(n24824), .O(n24825) );
  AOI22S U26352 ( .A1(n27685), .A2(img[198]), .B1(n29096), .B2(n30296), .O(
        n24826) );
  ND2S U26353 ( .I1(n25327), .I2(n24826), .O(n24827) );
  MUX2 U26354 ( .A(img[190]), .B(n24827), .S(n28848), .O(n13346) );
  AOI22S U26355 ( .A1(n26855), .A2(img[190]), .B1(n13781), .B2(n30297), .O(
        n24828) );
  ND2S U26356 ( .I1(n25327), .I2(n24828), .O(n24829) );
  MUX2 U26357 ( .A(img[198]), .B(n24829), .S(n28845), .O(n13334) );
  AOI22S U26358 ( .A1(n28347), .A2(img[326]), .B1(n28695), .B2(n30298), .O(
        n24830) );
  ND2S U26359 ( .I1(n25327), .I2(n24830), .O(n24831) );
  AOI22S U26360 ( .A1(n29435), .A2(img[318]), .B1(n28037), .B2(n30299), .O(
        n24832) );
  ND2S U26361 ( .I1(n25327), .I2(n24832), .O(n24833) );
  MUX2 U26362 ( .A(img[326]), .B(n24833), .S(n28851), .O(n13210) );
  AOI22S U26363 ( .A1(n28083), .A2(img[454]), .B1(n13779), .B2(n30300), .O(
        n24834) );
  ND2S U26364 ( .I1(n25327), .I2(n24834), .O(n24835) );
  AOI22S U26365 ( .A1(n25810), .A2(img[446]), .B1(n25062), .B2(n30301), .O(
        n24836) );
  ND2S U26366 ( .I1(n25327), .I2(n24836), .O(n24837) );
  MUX2 U26367 ( .A(img[454]), .B(n24837), .S(n28857), .O(n13078) );
  AOI22S U26368 ( .A1(n29076), .A2(img[1534]), .B1(n13779), .B2(n30302), .O(
        n24838) );
  ND2S U26369 ( .I1(n25327), .I2(n24838), .O(n24839) );
  BUF12CK U26370 ( .I(n25298), .O(n25327) );
  AOI22S U26371 ( .A1(n28938), .A2(n30303), .B1(n24890), .B2(img[1414]), .O(
        n24841) );
  ND3S U26372 ( .I1(n25327), .I2(n24841), .I3(n24840), .O(n24842) );
  MUX2 U26373 ( .A(img[1534]), .B(n24842), .S(n28868), .O(n12002) );
  AOI22S U26374 ( .A1(n27746), .A2(img[1478]), .B1(n23941), .B2(n30304), .O(
        n24843) );
  ND2S U26375 ( .I1(n25327), .I2(n24843), .O(n24844) );
  MUX2 U26376 ( .A(img[1470]), .B(n24844), .S(n28875), .O(n12066) );
  AOI22S U26377 ( .A1(n25062), .A2(n30305), .B1(n24890), .B2(img[1470]), .O(
        n24846) );
  ND3S U26378 ( .I1(n25327), .I2(n24846), .I3(n24845), .O(n24847) );
  MUX2 U26379 ( .A(img[1478]), .B(n24847), .S(n28872), .O(n12054) );
  INV1S U26380 ( .I(img[830]), .O(n24848) );
  AOI22S U26381 ( .A1(n26101), .A2(img[838]), .B1(n23941), .B2(n24848), .O(
        n24849) );
  ND2S U26382 ( .I1(n25327), .I2(n24849), .O(n24850) );
  MUX2 U26383 ( .A(n24850), .B(img[830]), .S(n28883), .O(n12702) );
  INV1S U26384 ( .I(img[838]), .O(n24851) );
  AOI22S U26385 ( .A1(n28347), .A2(img[830]), .B1(n24193), .B2(n24851), .O(
        n24852) );
  ND2S U26386 ( .I1(n25327), .I2(n24852), .O(n24853) );
  AOI22S U26387 ( .A1(n25595), .A2(img[710]), .B1(n23941), .B2(n30306), .O(
        n24854) );
  ND2S U26388 ( .I1(n25327), .I2(n24854), .O(n24855) );
  AOI22S U26389 ( .A1(n28083), .A2(img[702]), .B1(n13781), .B2(n30307), .O(
        n24856) );
  ND2S U26390 ( .I1(n25327), .I2(n24856), .O(n24857) );
  AOI22S U26391 ( .A1(n29129), .A2(img[1886]), .B1(n28695), .B2(n30308), .O(
        n24858) );
  ND2S U26392 ( .I1(n25327), .I2(n24858), .O(n24859) );
  MUX2 U26393 ( .A(n24859), .B(img[1830]), .S(n28892), .O(n11706) );
  AOI22S U26394 ( .A1(n27735), .A2(n30309), .B1(n24890), .B2(img[1830]), .O(
        n24861) );
  ND2S U26395 ( .I1(n13770), .I2(img[1894]), .O(n24860) );
  ND3S U26396 ( .I1(n25327), .I2(n24861), .I3(n24860), .O(n24862) );
  AOI22S U26397 ( .A1(n27990), .A2(img[1894]), .B1(n24193), .B2(n30310), .O(
        n24863) );
  ND2S U26398 ( .I1(n25327), .I2(n24863), .O(n24864) );
  AOI22S U26399 ( .A1(n29397), .A2(n30311), .B1(n24890), .B2(img[1822]), .O(
        n24866) );
  AOI22S U26400 ( .A1(n13901), .A2(img[1886]), .B1(img[1918]), .B2(n13782), 
        .O(n24865) );
  ND3S U26401 ( .I1(n25327), .I2(n24866), .I3(n24865), .O(n24867) );
  MUX2 U26402 ( .A(img[1894]), .B(n24867), .S(n28903), .O(n11642) );
  AOI22S U26403 ( .A1(n29435), .A2(img[1918]), .B1(n24374), .B2(n30312), .O(
        n24868) );
  ND2S U26404 ( .I1(n25327), .I2(n24868), .O(n24869) );
  MUX2 U26405 ( .A(img[1798]), .B(n24869), .S(n28906), .O(n11738) );
  AOI22S U26406 ( .A1(n27735), .A2(n30313), .B1(n24890), .B2(img[1798]), .O(
        n24871) );
  AOI22S U26407 ( .A1(n13899), .A2(img[1862]), .B1(img[1894]), .B2(n13782), 
        .O(n24870) );
  ND3S U26408 ( .I1(n25327), .I2(n24871), .I3(n24870), .O(n24872) );
  MUX2 U26409 ( .A(img[1918]), .B(n24872), .S(n28911), .O(n11614) );
  AOI22S U26410 ( .A1(n27685), .A2(img[1862]), .B1(n24374), .B2(n30314), .O(
        n24873) );
  ND2S U26411 ( .I1(n25327), .I2(n24873), .O(n24874) );
  MUX2 U26412 ( .A(img[1854]), .B(n24874), .S(n28919), .O(n11678) );
  AOI22S U26413 ( .A1(n29407), .A2(n30315), .B1(n24890), .B2(img[1854]), .O(
        n24876) );
  ND3S U26414 ( .I1(n25327), .I2(n24876), .I3(n24875), .O(n24877) );
  MUX2 U26415 ( .A(img[1862]), .B(n24877), .S(n28916), .O(n11674) );
  AOI22S U26416 ( .A1(n13773), .A2(img[1758]), .B1(n24193), .B2(n30316), .O(
        n24878) );
  ND2S U26417 ( .I1(n25327), .I2(n24878), .O(n24879) );
  MUX2 U26418 ( .A(n24879), .B(img[1702]), .S(n28922), .O(n11830) );
  AOI22S U26419 ( .A1(n28913), .A2(n30317), .B1(n24890), .B2(img[1702]), .O(
        n24881) );
  ND2S U26420 ( .I1(n13770), .I2(img[1766]), .O(n24880) );
  ND3S U26421 ( .I1(n25327), .I2(n24881), .I3(n24880), .O(n24882) );
  AOI22S U26422 ( .A1(n28347), .A2(img[1766]), .B1(n29096), .B2(n30318), .O(
        n24883) );
  ND2S U26423 ( .I1(n25327), .I2(n24883), .O(n24884) );
  AOI22S U26424 ( .A1(n25377), .A2(n30319), .B1(n24890), .B2(img[1694]), .O(
        n24886) );
  AOI22S U26425 ( .A1(n13903), .A2(img[1758]), .B1(img[1790]), .B2(n13782), 
        .O(n24885) );
  ND3S U26426 ( .I1(n25327), .I2(n24886), .I3(n24885), .O(n24887) );
  MUX2 U26427 ( .A(img[1766]), .B(n24887), .S(n28933), .O(n11766) );
  AOI22S U26428 ( .A1(n24415), .A2(img[1790]), .B1(n29397), .B2(n30320), .O(
        n24888) );
  ND2S U26429 ( .I1(n25327), .I2(n24888), .O(n24889) );
  AOI22S U26430 ( .A1(n25377), .A2(n30321), .B1(n24890), .B2(img[1670]), .O(
        n24892) );
  AOI22S U26431 ( .A1(n13904), .A2(img[1734]), .B1(img[1766]), .B2(n13782), 
        .O(n24891) );
  ND3S U26432 ( .I1(n25327), .I2(n24892), .I3(n24891), .O(n24893) );
  MUX2 U26433 ( .A(img[1790]), .B(n24893), .S(n28941), .O(n11746) );
  AOI22S U26434 ( .A1(n28347), .A2(img[1734]), .B1(n13781), .B2(n30322), .O(
        n24894) );
  ND2S U26435 ( .I1(n25327), .I2(n24894), .O(n24895) );
  AOI22S U26436 ( .A1(n29397), .A2(n30323), .B1(n24946), .B2(img[1726]), .O(
        n24897) );
  ND2S U26437 ( .I1(n13902), .I2(img[1790]), .O(n24896) );
  ND3S U26438 ( .I1(n25327), .I2(n24897), .I3(n24896), .O(n24898) );
  MUX2 U26439 ( .A(img[1734]), .B(n24898), .S(n28945), .O(n11798) );
  AOI22S U26440 ( .A1(n29076), .A2(img[1630]), .B1(n13781), .B2(n30324), .O(
        n24899) );
  ND2S U26441 ( .I1(n25327), .I2(n24899), .O(n24900) );
  MUX2 U26442 ( .A(n24900), .B(img[1574]), .S(n28951), .O(n11962) );
  AOI22S U26443 ( .A1(n29242), .A2(n30325), .B1(n24946), .B2(img[1574]), .O(
        n24902) );
  ND3S U26444 ( .I1(n25327), .I2(n24902), .I3(n24901), .O(n24903) );
  AOI22S U26445 ( .A1(n25595), .A2(img[1638]), .B1(n13781), .B2(n30326), .O(
        n24904) );
  ND2S U26446 ( .I1(n25327), .I2(n24904), .O(n24905) );
  AOI22S U26447 ( .A1(n29242), .A2(n30327), .B1(n24946), .B2(img[1566]), .O(
        n24907) );
  AOI22S U26448 ( .A1(n13905), .A2(img[1630]), .B1(img[1662]), .B2(n13782), 
        .O(n24906) );
  ND3S U26449 ( .I1(n25327), .I2(n24907), .I3(n24906), .O(n24908) );
  MUX2 U26450 ( .A(img[1638]), .B(n24908), .S(n28962), .O(n11897) );
  AOI22S U26451 ( .A1(n25595), .A2(img[1662]), .B1(n13781), .B2(n30328), .O(
        n24909) );
  ND2S U26452 ( .I1(n25327), .I2(n24909), .O(n24910) );
  AOI22S U26453 ( .A1(n29242), .A2(n30329), .B1(n24946), .B2(img[1542]), .O(
        n24912) );
  AOI22S U26454 ( .A1(n13903), .A2(img[1606]), .B1(img[1638]), .B2(n28908), 
        .O(n24911) );
  ND3S U26455 ( .I1(n25327), .I2(n24912), .I3(n24911), .O(n24913) );
  MUX2 U26456 ( .A(img[1662]), .B(n24913), .S(n28969), .O(n11870) );
  AOI22S U26457 ( .A1(n13777), .A2(img[1606]), .B1(n13781), .B2(n30330), .O(
        n24914) );
  ND2S U26458 ( .I1(n25327), .I2(n24914), .O(n24915) );
  MUX2 U26459 ( .A(img[1598]), .B(n24915), .S(n28976), .O(n11934) );
  AOI22S U26460 ( .A1(n28695), .A2(n30331), .B1(n24946), .B2(img[1598]), .O(
        n24917) );
  ND3S U26461 ( .I1(n25327), .I2(n24917), .I3(n24916), .O(n24918) );
  MUX2 U26462 ( .A(img[1606]), .B(n24918), .S(n28973), .O(n11930) );
  AOI22S U26463 ( .A1(n13776), .A2(img[1150]), .B1(n27735), .B2(n30332), .O(
        n24919) );
  ND2S U26464 ( .I1(n25327), .I2(n24919), .O(n24920) );
  AOI22S U26465 ( .A1(n28695), .A2(n30333), .B1(n24946), .B2(img[1030]), .O(
        n24922) );
  ND3S U26466 ( .I1(n25327), .I2(n24922), .I3(n24921), .O(n24923) );
  MUX2 U26467 ( .A(img[1150]), .B(n24923), .S(n28983), .O(n12382) );
  AOI22S U26468 ( .A1(n27957), .A2(img[1094]), .B1(n28075), .B2(n30334), .O(
        n24924) );
  ND2S U26469 ( .I1(n25327), .I2(n24924), .O(n24925) );
  MUX2 U26470 ( .A(img[1086]), .B(n24925), .S(n28990), .O(n12446) );
  AOI22S U26471 ( .A1(n28695), .A2(n30335), .B1(n24946), .B2(img[1086]), .O(
        n24927) );
  ND3S U26472 ( .I1(n25327), .I2(n24927), .I3(n24926), .O(n24928) );
  MUX2 U26473 ( .A(img[1094]), .B(n24928), .S(n28987), .O(n12439) );
  AOI22S U26474 ( .A1(n26855), .A2(img[2014]), .B1(n28162), .B2(n30336), .O(
        n24929) );
  ND2S U26475 ( .I1(n25327), .I2(n24929), .O(n24930) );
  MUX2 U26476 ( .A(n24930), .B(img[1958]), .S(n28993), .O(n11574) );
  AOI22S U26477 ( .A1(n28695), .A2(n30337), .B1(n24946), .B2(img[1958]), .O(
        n24932) );
  ND3S U26478 ( .I1(n25327), .I2(n24932), .I3(n24931), .O(n24933) );
  AOI22S U26479 ( .A1(n26101), .A2(img[2022]), .B1(n29242), .B2(n30338), .O(
        n24934) );
  ND2S U26480 ( .I1(n25327), .I2(n24934), .O(n24935) );
  MUX2 U26481 ( .A(img[1950]), .B(n24935), .S(n29000), .O(n11586) );
  AOI22S U26482 ( .A1(n28695), .A2(n30339), .B1(n24946), .B2(img[1950]), .O(
        n24937) );
  AOI22S U26483 ( .A1(n13899), .A2(img[2014]), .B1(img[2046]), .B2(n13782), 
        .O(n24936) );
  ND3S U26484 ( .I1(n25327), .I2(n24937), .I3(n24936), .O(n24938) );
  MUX2 U26485 ( .A(img[2022]), .B(n24938), .S(n29004), .O(n11510) );
  AOI22S U26486 ( .A1(n28347), .A2(img[2046]), .B1(n13781), .B2(n30340), .O(
        n24939) );
  ND2S U26487 ( .I1(n25327), .I2(n24939), .O(n24940) );
  MUX2 U26488 ( .A(img[1926]), .B(n24940), .S(n29007), .O(n11606) );
  AOI22S U26489 ( .A1(n28695), .A2(n30341), .B1(n24946), .B2(img[1926]), .O(
        n24942) );
  AOI22S U26490 ( .A1(n13903), .A2(img[1990]), .B1(img[2022]), .B2(n13782), 
        .O(n24941) );
  ND3S U26491 ( .I1(n25327), .I2(n24942), .I3(n24941), .O(n24943) );
  AOI22S U26492 ( .A1(n28643), .A2(img[1990]), .B1(n13781), .B2(n30342), .O(
        n24944) );
  ND2S U26493 ( .I1(n25327), .I2(n24944), .O(n24945) );
  MUX2 U26494 ( .A(img[1982]), .B(n24945), .S(n29018), .O(n11554) );
  AOI22S U26495 ( .A1(n28695), .A2(n30343), .B1(n24946), .B2(img[1982]), .O(
        n24948) );
  ND2S U26496 ( .I1(n29124), .I2(img[2046]), .O(n24947) );
  ND3S U26497 ( .I1(n25327), .I2(n24948), .I3(n24947), .O(n24949) );
  MUX2 U26498 ( .A(img[1990]), .B(n24949), .S(n29015), .O(n11542) );
  AOI22S U26499 ( .A1(n27722), .A2(img[630]), .B1(n29242), .B2(n30344), .O(
        n24950) );
  ND2S U26500 ( .I1(n25327), .I2(n24950), .O(n24951) );
  AOI22S U26501 ( .A1(n27746), .A2(img[526]), .B1(n25859), .B2(n30345), .O(
        n24952) );
  ND2S U26502 ( .I1(n25327), .I2(n24952), .O(n24953) );
  MUX2 U26503 ( .A(n24953), .B(img[630]), .S(n29292), .O(n12906) );
  AOI22S U26504 ( .A1(n28347), .A2(img[118]), .B1(n29397), .B2(n30346), .O(
        n24954) );
  ND2S U26505 ( .I1(n25327), .I2(n24954), .O(n24955) );
  AOI22S U26506 ( .A1(n26855), .A2(img[14]), .B1(n27511), .B2(n30347), .O(
        n24956) );
  ND2S U26507 ( .I1(n25327), .I2(n24956), .O(n24959) );
  MUX2 U26508 ( .A(img[118]), .B(n24959), .S(n29536), .O(n13418) );
  AOI22S U26509 ( .A1(n13771), .A2(img[1230]), .B1(n13781), .B2(n30348), .O(
        n24960) );
  ND2S U26510 ( .I1(n25327), .I2(n24960), .O(n24961) );
  AOI22S U26511 ( .A1(n25591), .A2(n30349), .B1(n24313), .B2(img[1206]), .O(
        n24963) );
  ND2S U26512 ( .I1(n29124), .I2(img[1270]), .O(n24962) );
  ND3S U26513 ( .I1(n25327), .I2(n24963), .I3(n24962), .O(n24964) );
  MUX2 U26514 ( .A(img[1230]), .B(n24964), .S(n28602), .O(n12306) );
  AOI22S U26515 ( .A1(n26855), .A2(img[1270]), .B1(n27511), .B2(n30350), .O(
        n24965) );
  ND2S U26516 ( .I1(n25327), .I2(n24965), .O(n24966) );
  AOI22S U26517 ( .A1(n25591), .A2(n30351), .B1(n25444), .B2(img[1166]), .O(
        n24968) );
  ND2S U26518 ( .I1(n29124), .I2(img[1230]), .O(n24967) );
  ND3S U26519 ( .I1(n25327), .I2(n24968), .I3(n24967), .O(n24969) );
  MUX2 U26520 ( .A(img[1270]), .B(n24969), .S(n28595), .O(n12262) );
  AOI22S U26521 ( .A1(n13773), .A2(img[1358]), .B1(n28862), .B2(n30352), .O(
        n24970) );
  ND2S U26522 ( .I1(n25327), .I2(n24970), .O(n24971) );
  MUX2 U26523 ( .A(n24971), .B(img[1334]), .S(n28612), .O(n12202) );
  AOI22S U26524 ( .A1(n25591), .A2(n30353), .B1(n25444), .B2(img[1334]), .O(
        n24973) );
  ND2S U26525 ( .I1(n29124), .I2(img[1398]), .O(n24972) );
  ND3S U26526 ( .I1(n25327), .I2(n24973), .I3(n24972), .O(n24974) );
  MUX2 U26527 ( .A(img[1358]), .B(n24974), .S(n28617), .O(n12174) );
  AOI22S U26528 ( .A1(n27065), .A2(img[1398]), .B1(n28913), .B2(n30354), .O(
        n24975) );
  ND2S U26529 ( .I1(n25327), .I2(n24975), .O(n24976) );
  AOI22S U26530 ( .A1(n25591), .A2(n30355), .B1(n28069), .B2(img[1294]), .O(
        n24978) );
  ND2S U26531 ( .I1(n29124), .I2(img[1358]), .O(n24977) );
  ND3S U26532 ( .I1(n25327), .I2(n24978), .I3(n24977), .O(n24979) );
  MUX2 U26533 ( .A(img[1398]), .B(n24979), .S(n28609), .O(n12138) );
  AOI22S U26534 ( .A1(n25810), .A2(img[1014]), .B1(n24193), .B2(n30356), .O(
        n24980) );
  ND2S U26535 ( .I1(n25327), .I2(n24980), .O(n24981) );
  MUX2 U26536 ( .A(img[910]), .B(n24981), .S(n29300), .O(n12626) );
  AOI22S U26537 ( .A1(n24415), .A2(img[910]), .B1(n13781), .B2(n30357), .O(
        n24982) );
  ND2S U26538 ( .I1(n25327), .I2(n24982), .O(n24983) );
  AOI22S U26539 ( .A1(n25810), .A2(img[246]), .B1(n13781), .B2(n30358), .O(
        n24984) );
  ND2S U26540 ( .I1(n25327), .I2(n24984), .O(n24985) );
  AOI22S U26541 ( .A1(n29414), .A2(img[142]), .B1(n13781), .B2(n30359), .O(
        n24986) );
  ND2S U26542 ( .I1(n25327), .I2(n24986), .O(n24987) );
  MUX2 U26543 ( .A(img[246]), .B(n24987), .S(n29309), .O(n13286) );
  AOI22S U26544 ( .A1(n26970), .A2(img[374]), .B1(n28913), .B2(n30360), .O(
        n24988) );
  ND2S U26545 ( .I1(n25327), .I2(n24988), .O(n24989) );
  MUX2 U26546 ( .A(n24989), .B(img[270]), .S(n29312), .O(n13262) );
  AOI22S U26547 ( .A1(n26101), .A2(img[270]), .B1(n13779), .B2(n30361), .O(
        n24990) );
  ND2S U26548 ( .I1(n25327), .I2(n24990), .O(n24991) );
  AOI22S U26549 ( .A1(n24415), .A2(img[502]), .B1(n28862), .B2(n30362), .O(
        n24992) );
  ND2S U26550 ( .I1(n25327), .I2(n24992), .O(n24993) );
  MUX2 U26551 ( .A(n24993), .B(img[398]), .S(n29318), .O(n13138) );
  AOI22S U26552 ( .A1(n28840), .A2(img[398]), .B1(n29457), .B2(n30363), .O(
        n24994) );
  ND2S U26553 ( .I1(n25327), .I2(n24994), .O(n24995) );
  MUX2 U26554 ( .A(img[502]), .B(n24995), .S(n29321), .O(n13030) );
  AOI22S U26555 ( .A1(n28840), .A2(img[1486]), .B1(n28862), .B2(n30364), .O(
        n24996) );
  ND2S U26556 ( .I1(n25327), .I2(n24996), .O(n24997) );
  AOI22S U26557 ( .A1(n28614), .A2(n30365), .B1(n28043), .B2(img[1462]), .O(
        n24999) );
  ND2S U26558 ( .I1(n29124), .I2(img[1526]), .O(n24998) );
  ND3S U26559 ( .I1(n25327), .I2(n24999), .I3(n24998), .O(n25000) );
  MUX2 U26560 ( .A(img[1486]), .B(n25000), .S(n28656), .O(n12050) );
  AOI22S U26561 ( .A1(n26822), .A2(img[1526]), .B1(n28913), .B2(n30366), .O(
        n25001) );
  ND2S U26562 ( .I1(n25327), .I2(n25001), .O(n25002) );
  MUX2 U26563 ( .A(n25002), .B(img[1422]), .S(n28645), .O(n12114) );
  AOI22S U26564 ( .A1(n28614), .A2(n30367), .B1(n28069), .B2(img[1422]), .O(
        n25004) );
  ND3S U26565 ( .I1(n25327), .I2(n25004), .I3(n25003), .O(n25005) );
  AOI22S U26566 ( .A1(n26822), .A2(img[886]), .B1(n29457), .B2(n30368), .O(
        n25006) );
  ND2S U26567 ( .I1(n25327), .I2(n25006), .O(n25007) );
  MUX2 U26568 ( .A(img[782]), .B(n25007), .S(n29324), .O(n12750) );
  INV1S U26569 ( .I(img[886]), .O(n25008) );
  AOI22S U26570 ( .A1(n28382), .A2(img[782]), .B1(n13779), .B2(n25008), .O(
        n25009) );
  ND2S U26571 ( .I1(n25327), .I2(n25009), .O(n25010) );
  AOI22S U26572 ( .A1(n28083), .A2(img[758]), .B1(n13779), .B2(n30369), .O(
        n25011) );
  ND2S U26573 ( .I1(n25327), .I2(n25011), .O(n25012) );
  AOI22S U26574 ( .A1(n28318), .A2(img[654]), .B1(n29407), .B2(n30370), .O(
        n25013) );
  ND2S U26575 ( .I1(n25327), .I2(n25013), .O(n25014) );
  AOI22S U26576 ( .A1(n13776), .A2(img[1878]), .B1(n25377), .B2(n30371), .O(
        n25015) );
  ND2S U26577 ( .I1(n25327), .I2(n25015), .O(n25016) );
  MUX2 U26578 ( .A(n25016), .B(img[1838]), .S(n28672), .O(n11694) );
  AOI22S U26579 ( .A1(n25591), .A2(n30372), .B1(n24434), .B2(img[1838]), .O(
        n25018) );
  ND2S U26580 ( .I1(n29124), .I2(img[1902]), .O(n25017) );
  ND3S U26581 ( .I1(n25327), .I2(n25018), .I3(n25017), .O(n25019) );
  MUX2 U26582 ( .A(img[1878]), .B(n25019), .S(n28676), .O(n11658) );
  AOI22S U26583 ( .A1(n13780), .A2(img[1902]), .B1(n28162), .B2(n30373), .O(
        n25020) );
  ND2S U26584 ( .I1(n25327), .I2(n25020), .O(n25021) );
  MUX2 U26585 ( .A(n25021), .B(img[1814]), .S(n28679), .O(n11722) );
  AOI22S U26586 ( .A1(n29194), .A2(n30374), .B1(n28069), .B2(img[1814]), .O(
        n25023) );
  AOI22S U26587 ( .A1(n13904), .A2(img[1878]), .B1(img[1910]), .B2(n13782), 
        .O(n25022) );
  ND3S U26588 ( .I1(n25327), .I2(n25023), .I3(n25022), .O(n25024) );
  MUX2 U26589 ( .A(img[1902]), .B(n25024), .S(n28683), .O(n11630) );
  AOI22S U26590 ( .A1(n13780), .A2(img[1870]), .B1(n28037), .B2(n30375), .O(
        n25025) );
  ND2S U26591 ( .I1(n25168), .I2(n25025), .O(n25026) );
  MUX2 U26592 ( .A(n25026), .B(img[1846]), .S(n28693), .O(n11690) );
  AOI22S U26593 ( .A1(n25062), .A2(n30376), .B1(n24313), .B2(img[1846]), .O(
        n25028) );
  ND3S U26594 ( .I1(n25327), .I2(n25028), .I3(n25027), .O(n25029) );
  MUX2 U26595 ( .A(img[1870]), .B(n25029), .S(n28698), .O(n11662) );
  AOI22S U26596 ( .A1(n26970), .A2(img[1910]), .B1(n28075), .B2(n30377), .O(
        n25030) );
  ND2S U26597 ( .I1(n25327), .I2(n25030), .O(n25031) );
  AOI22S U26598 ( .A1(n28592), .A2(n30378), .B1(n28069), .B2(img[1806]), .O(
        n25033) );
  AOI22S U26599 ( .A1(n13903), .A2(img[1870]), .B1(img[1902]), .B2(n13782), 
        .O(n25032) );
  ND3S U26600 ( .I1(n25327), .I2(n25033), .I3(n25032), .O(n25034) );
  MUX2 U26601 ( .A(img[1910]), .B(n25034), .S(n28690), .O(n11626) );
  AOI22S U26602 ( .A1(n26101), .A2(img[1750]), .B1(n28075), .B2(n30379), .O(
        n25035) );
  ND2S U26603 ( .I1(n25327), .I2(n25035), .O(n25036) );
  AOI22S U26604 ( .A1(n28592), .A2(n30380), .B1(n28069), .B2(img[1710]), .O(
        n25038) );
  ND2S U26605 ( .I1(n29124), .I2(img[1774]), .O(n25037) );
  ND3S U26606 ( .I1(n25327), .I2(n25038), .I3(n25037), .O(n25039) );
  MUX2 U26607 ( .A(img[1750]), .B(n25039), .S(n28705), .O(n11782) );
  AOI22S U26608 ( .A1(n28347), .A2(img[1774]), .B1(n28075), .B2(n30381), .O(
        n25040) );
  ND2S U26609 ( .I1(n25327), .I2(n25040), .O(n25041) );
  AOI22S U26610 ( .A1(n28592), .A2(n30382), .B1(n29257), .B2(img[1686]), .O(
        n25043) );
  AOI22S U26611 ( .A1(n13770), .A2(img[1750]), .B1(img[1782]), .B2(n13782), 
        .O(n25042) );
  ND3S U26612 ( .I1(n25327), .I2(n25043), .I3(n25042), .O(n25044) );
  MUX2 U26613 ( .A(img[1774]), .B(n25044), .S(n28712), .O(n11762) );
  AOI22S U26614 ( .A1(n25595), .A2(img[1742]), .B1(n28075), .B2(n30383), .O(
        n25045) );
  ND2S U26615 ( .I1(n25327), .I2(n25045), .O(n25046) );
  MUX2 U26616 ( .A(n25046), .B(img[1718]), .S(n28722), .O(n11814) );
  AOI22S U26617 ( .A1(n28592), .A2(n30384), .B1(n24808), .B2(img[1718]), .O(
        n25048) );
  ND2S U26618 ( .I1(n29124), .I2(img[1782]), .O(n25047) );
  ND3S U26619 ( .I1(n25327), .I2(n25048), .I3(n25047), .O(n25049) );
  MUX2 U26620 ( .A(img[1742]), .B(n25049), .S(n28726), .O(n11794) );
  AOI22S U26621 ( .A1(n29435), .A2(img[1782]), .B1(n28075), .B2(n30385), .O(
        n25050) );
  ND2S U26622 ( .I1(n25327), .I2(n25050), .O(n25051) );
  AOI22S U26623 ( .A1(n28592), .A2(n30386), .B1(n24946), .B2(img[1678]), .O(
        n25053) );
  AOI22S U26624 ( .A1(n13905), .A2(img[1742]), .B1(img[1774]), .B2(n13782), 
        .O(n25052) );
  ND3S U26625 ( .I1(n25327), .I2(n25053), .I3(n25052), .O(n25054) );
  MUX2 U26626 ( .A(img[1782]), .B(n25054), .S(n28719), .O(n11750) );
  AOI22S U26627 ( .A1(n29072), .A2(img[1622]), .B1(n28037), .B2(n30387), .O(
        n25055) );
  ND2S U26628 ( .I1(n25327), .I2(n25055), .O(n25056) );
  MUX2 U26629 ( .A(n25056), .B(img[1582]), .S(n28729), .O(n11950) );
  AOI22S U26630 ( .A1(n28592), .A2(n30388), .B1(n28069), .B2(img[1582]), .O(
        n25058) );
  ND3S U26631 ( .I1(n25327), .I2(n25058), .I3(n25057), .O(n25059) );
  MUX2 U26632 ( .A(img[1622]), .B(n25059), .S(n28733), .O(n11914) );
  AOI22S U26633 ( .A1(n28412), .A2(img[1646]), .B1(n28037), .B2(n30389), .O(
        n25060) );
  ND2S U26634 ( .I1(n25327), .I2(n25060), .O(n25061) );
  MUX2 U26635 ( .A(n25061), .B(img[1558]), .S(n28736), .O(n11978) );
  AOI22S U26636 ( .A1(n28938), .A2(n30390), .B1(n24946), .B2(img[1558]), .O(
        n25064) );
  AOI22S U26637 ( .A1(n13903), .A2(img[1622]), .B1(img[1654]), .B2(n13782), 
        .O(n25063) );
  ND3S U26638 ( .I1(n25327), .I2(n25064), .I3(n25063), .O(n25065) );
  MUX2 U26639 ( .A(img[1646]), .B(n25065), .S(n28740), .O(n11886) );
  AOI22S U26640 ( .A1(n27065), .A2(img[1614]), .B1(n28037), .B2(n30391), .O(
        n25066) );
  ND2S U26641 ( .I1(n25327), .I2(n25066), .O(n25067) );
  AOI22S U26642 ( .A1(n25062), .A2(n30392), .B1(n26091), .B2(img[1590]), .O(
        n25069) );
  ND2S U26643 ( .I1(n29124), .I2(img[1654]), .O(n25068) );
  ND3 U26644 ( .I1(n25298), .I2(n25069), .I3(n25068), .O(n25070) );
  AOI22S U26645 ( .A1(n25595), .A2(img[1654]), .B1(n13781), .B2(n30393), .O(
        n25071) );
  ND2S U26646 ( .I1(n25327), .I2(n25071), .O(n25072) );
  AOI22S U26647 ( .A1(n25062), .A2(n30394), .B1(n28043), .B2(img[1550]), .O(
        n25074) );
  AOI22S U26648 ( .A1(n13904), .A2(img[1614]), .B1(img[1646]), .B2(n13782), 
        .O(n25073) );
  ND3S U26649 ( .I1(n25327), .I2(n25074), .I3(n25073), .O(n25075) );
  MUX2 U26650 ( .A(img[1654]), .B(n25075), .S(n28747), .O(n11882) );
  AOI22S U26651 ( .A1(n29072), .A2(img[1102]), .B1(n13775), .B2(n30395), .O(
        n25076) );
  ND2S U26652 ( .I1(n25327), .I2(n25076), .O(n25077) );
  MUX2 U26653 ( .A(n25077), .B(img[1078]), .S(n28764), .O(n12458) );
  AOI22S U26654 ( .A1(n25062), .A2(n30396), .B1(n24313), .B2(img[1078]), .O(
        n25079) );
  ND3S U26655 ( .I1(n25327), .I2(n25079), .I3(n25078), .O(n25080) );
  MUX2 U26656 ( .A(img[1102]), .B(n25080), .S(n28768), .O(n12430) );
  AOI22S U26657 ( .A1(n28643), .A2(img[1142]), .B1(n29407), .B2(n30397), .O(
        n25081) );
  ND2S U26658 ( .I1(n25327), .I2(n25081), .O(n25082) );
  AOI22S U26659 ( .A1(n25062), .A2(n30398), .B1(n24313), .B2(img[1038]), .O(
        n25084) );
  ND3S U26660 ( .I1(n25327), .I2(n25084), .I3(n25083), .O(n25085) );
  MUX2 U26661 ( .A(img[1142]), .B(n25085), .S(n28761), .O(n12394) );
  AOI22S U26662 ( .A1(n13777), .A2(img[2006]), .B1(n25591), .B2(n30399), .O(
        n25086) );
  ND2S U26663 ( .I1(n25327), .I2(n25086), .O(n25087) );
  MUX2 U26664 ( .A(n25087), .B(img[1966]), .S(n28771), .O(n11570) );
  AOI22S U26665 ( .A1(n25062), .A2(n30400), .B1(n24313), .B2(img[1966]), .O(
        n25089) );
  ND3S U26666 ( .I1(n25327), .I2(n25089), .I3(n25088), .O(n25090) );
  MUX2 U26667 ( .A(img[2006]), .B(n25090), .S(n28775), .O(n11526) );
  AOI22S U26668 ( .A1(n28083), .A2(img[2030]), .B1(n28075), .B2(n30401), .O(
        n25091) );
  ND2S U26669 ( .I1(n25327), .I2(n25091), .O(n25092) );
  MUX2 U26670 ( .A(n25092), .B(img[1942]), .S(n28778), .O(n11590) );
  AOI22S U26671 ( .A1(n25062), .A2(n30402), .B1(n28069), .B2(img[1942]), .O(
        n25094) );
  AOI22S U26672 ( .A1(n13899), .A2(img[2006]), .B1(img[2038]), .B2(n13782), 
        .O(n25093) );
  ND3S U26673 ( .I1(n25327), .I2(n25094), .I3(n25093), .O(n25095) );
  MUX2 U26674 ( .A(img[2030]), .B(n25095), .S(n28782), .O(n11506) );
  AOI22S U26675 ( .A1(n13778), .A2(img[1998]), .B1(n13781), .B2(n30403), .O(
        n25096) );
  ND2S U26676 ( .I1(n25327), .I2(n25096), .O(n25097) );
  MUX2 U26677 ( .A(n25097), .B(img[1974]), .S(n28792), .O(n11558) );
  AOI22S U26678 ( .A1(n27443), .A2(n30404), .B1(n24946), .B2(img[1974]), .O(
        n25099) );
  ND3S U26679 ( .I1(n25327), .I2(n25099), .I3(n25098), .O(n25100) );
  MUX2 U26680 ( .A(img[1998]), .B(n25100), .S(n28796), .O(n11538) );
  AOI22S U26681 ( .A1(n29435), .A2(img[2038]), .B1(n28433), .B2(n30405), .O(
        n25101) );
  ND2S U26682 ( .I1(n25168), .I2(n25101), .O(n25102) );
  MUX2 U26683 ( .A(img[1934]), .B(n25102), .S(n28785), .O(n11602) );
  AOI22S U26684 ( .A1(n27443), .A2(n30406), .B1(n24946), .B2(img[1934]), .O(
        n25104) );
  AOI22S U26685 ( .A1(n13899), .A2(img[1998]), .B1(img[2030]), .B2(n13782), 
        .O(n25103) );
  ND3S U26686 ( .I1(n25327), .I2(n25104), .I3(n25103), .O(n25105) );
  MUX2 U26687 ( .A(img[2038]), .B(n25105), .S(n28789), .O(n11494) );
  AOI22S U26688 ( .A1(n27110), .A2(img[542]), .B1(n28182), .B2(n30407), .O(
        n25106) );
  ND2S U26689 ( .I1(n25168), .I2(n25106), .O(n25107) );
  MUX2 U26690 ( .A(n25107), .B(img[614]), .S(n29286), .O(n12922) );
  BUF2 U26691 ( .I(n25298), .O(n25168) );
  AOI22S U26692 ( .A1(n28221), .A2(img[614]), .B1(n24755), .B2(n30408), .O(
        n25108) );
  ND2S U26693 ( .I1(n25168), .I2(n25108), .O(n25109) );
  AOI22S U26694 ( .A1(n26822), .A2(img[30]), .B1(n13781), .B2(n30409), .O(
        n25110) );
  ND2S U26695 ( .I1(n25168), .I2(n25110), .O(n25111) );
  MUX2 U26696 ( .A(img[102]), .B(n25111), .S(n29280), .O(n13434) );
  AOI22S U26697 ( .A1(n28318), .A2(img[102]), .B1(n13781), .B2(n30410), .O(
        n25112) );
  ND2S U26698 ( .I1(n25168), .I2(n25112), .O(n25113) );
  AOI22S U26699 ( .A1(n28347), .A2(img[1246]), .B1(n25062), .B2(n30411), .O(
        n25114) );
  ND2S U26700 ( .I1(n25168), .I2(n25114), .O(n25115) );
  MUX2 U26701 ( .A(n25115), .B(img[1190]), .S(n29207), .O(n12342) );
  AOI22S U26702 ( .A1(n27443), .A2(n30412), .B1(n28069), .B2(img[1190]), .O(
        n25117) );
  ND3S U26703 ( .I1(n25327), .I2(n25117), .I3(n25116), .O(n25118) );
  MUX2 U26704 ( .A(img[1246]), .B(n25118), .S(n29211), .O(n12290) );
  AOI22S U26705 ( .A1(n27443), .A2(n30413), .B1(n25444), .B2(img[1182]), .O(
        n25120) );
  ND3S U26706 ( .I1(n25327), .I2(n25120), .I3(n25119), .O(n25121) );
  MUX2 U26707 ( .A(img[1254]), .B(n25121), .S(n29218), .O(n12278) );
  AOI22S U26708 ( .A1(n27065), .A2(img[1254]), .B1(n25062), .B2(n30414), .O(
        n25122) );
  ND2S U26709 ( .I1(n25168), .I2(n25122), .O(n25123) );
  MUX2 U26710 ( .A(img[1182]), .B(n25123), .S(n29214), .O(n12354) );
  AOI22S U26711 ( .A1(n26970), .A2(img[1374]), .B1(n28037), .B2(n30415), .O(
        n25124) );
  ND2S U26712 ( .I1(n25168), .I2(n25124), .O(n25125) );
  MUX2 U26713 ( .A(n25125), .B(img[1318]), .S(n29233), .O(n12218) );
  AOI22S U26714 ( .A1(n27443), .A2(n30416), .B1(n25444), .B2(img[1318]), .O(
        n25127) );
  ND3S U26715 ( .I1(n25327), .I2(n25127), .I3(n25126), .O(n25128) );
  MUX2 U26716 ( .A(img[1374]), .B(n25128), .S(n29237), .O(n12158) );
  AOI22S U26717 ( .A1(n27443), .A2(n30417), .B1(n27919), .B2(img[1310]), .O(
        n25130) );
  ND3S U26718 ( .I1(n25327), .I2(n25130), .I3(n25129), .O(n25131) );
  MUX2 U26719 ( .A(img[1382]), .B(n25131), .S(n29245), .O(n12154) );
  AOI22S U26720 ( .A1(n28412), .A2(img[1382]), .B1(n27735), .B2(n30418), .O(
        n25132) );
  ND2S U26721 ( .I1(n25168), .I2(n25132), .O(n25133) );
  MUX2 U26722 ( .A(img[1310]), .B(n25133), .S(n29240), .O(n12222) );
  AOI22S U26723 ( .A1(n28412), .A2(img[926]), .B1(n27735), .B2(n30419), .O(
        n25134) );
  ND2S U26724 ( .I1(n25168), .I2(n25134), .O(n25135) );
  MUX2 U26725 ( .A(img[998]), .B(n25135), .S(n29224), .O(n12534) );
  AOI22S U26726 ( .A1(n28643), .A2(img[998]), .B1(n27735), .B2(n30420), .O(
        n25136) );
  ND2S U26727 ( .I1(n25168), .I2(n25136), .O(n25137) );
  AOI22S U26728 ( .A1(n28643), .A2(img[158]), .B1(n27735), .B2(n30421), .O(
        n25138) );
  ND2S U26729 ( .I1(n25168), .I2(n25138), .O(n25139) );
  MUX2 U26730 ( .A(img[230]), .B(n25139), .S(n29267), .O(n13302) );
  AOI22S U26731 ( .A1(n28643), .A2(img[230]), .B1(n27735), .B2(n30422), .O(
        n25140) );
  ND2S U26732 ( .I1(n25168), .I2(n25140), .O(n25141) );
  MUX2 U26733 ( .A(img[158]), .B(n25141), .S(n29264), .O(n13378) );
  AOI22S U26734 ( .A1(n28643), .A2(img[286]), .B1(n27735), .B2(n30423), .O(
        n25142) );
  ND2S U26735 ( .I1(n25168), .I2(n25142), .O(n25143) );
  MUX2 U26736 ( .A(img[358]), .B(n25143), .S(n29182), .O(n13178) );
  AOI22S U26737 ( .A1(n28643), .A2(img[358]), .B1(n27511), .B2(n30424), .O(
        n25144) );
  ND2S U26738 ( .I1(n25168), .I2(n25144), .O(n25145) );
  AOI22S U26739 ( .A1(n28643), .A2(img[414]), .B1(n23941), .B2(n30425), .O(
        n25146) );
  ND2S U26740 ( .I1(n25168), .I2(n25146), .O(n25147) );
  MUX2 U26741 ( .A(img[486]), .B(n25147), .S(n29273), .O(n13046) );
  AOI22S U26742 ( .A1(n28643), .A2(img[486]), .B1(n13781), .B2(n30426), .O(
        n25148) );
  ND2S U26743 ( .I1(n25168), .I2(n25148), .O(n25149) );
  AOI22S U26744 ( .A1(n24415), .A2(img[1502]), .B1(n23941), .B2(n30427), .O(
        n25150) );
  ND2S U26745 ( .I1(n25168), .I2(n25150), .O(n25151) );
  MUX2 U26746 ( .A(n25151), .B(img[1446]), .S(n29248), .O(n12086) );
  AOI22S U26747 ( .A1(n28135), .A2(n30428), .B1(n25444), .B2(img[1446]), .O(
        n25153) );
  ND3S U26748 ( .I1(n25327), .I2(n25153), .I3(n25152), .O(n25154) );
  AOI22S U26749 ( .A1(n28135), .A2(n30429), .B1(n27919), .B2(img[1438]), .O(
        n25156) );
  ND3S U26750 ( .I1(n25327), .I2(n25156), .I3(n25155), .O(n25157) );
  MUX2 U26751 ( .A(img[1510]), .B(n25157), .S(n29261), .O(n12022) );
  AOI22S U26752 ( .A1(n28840), .A2(img[1510]), .B1(n27735), .B2(n30430), .O(
        n25158) );
  ND2S U26753 ( .I1(n25168), .I2(n25158), .O(n25159) );
  MUX2 U26754 ( .A(n25159), .B(img[1438]), .S(n29255), .O(n12098) );
  INV1S U26755 ( .I(img[870]), .O(n25160) );
  AOI22S U26756 ( .A1(n29435), .A2(img[798]), .B1(n29194), .B2(n25160), .O(
        n25161) );
  ND2S U26757 ( .I1(n25168), .I2(n25161), .O(n25162) );
  AOI22S U26758 ( .A1(n28347), .A2(img[870]), .B1(n29194), .B2(n30431), .O(
        n25163) );
  ND2S U26759 ( .I1(n25168), .I2(n25163), .O(n25164) );
  MUX2 U26760 ( .A(img[798]), .B(n25164), .S(n29227), .O(n12734) );
  AOI22S U26761 ( .A1(n29072), .A2(img[670]), .B1(n25591), .B2(n30432), .O(
        n25165) );
  ND2S U26762 ( .I1(n25168), .I2(n25165), .O(n25166) );
  MUX2 U26763 ( .A(n25166), .B(img[742]), .S(n29204), .O(n12790) );
  AOI22S U26764 ( .A1(n28347), .A2(img[742]), .B1(n29530), .B2(n30433), .O(
        n25167) );
  ND2S U26765 ( .I1(n25168), .I2(n25167), .O(n25169) );
  BUF2 U26766 ( .I(n25298), .O(n25258) );
  AOI22S U26767 ( .A1(n28347), .A2(img[1118]), .B1(n29457), .B2(n30434), .O(
        n25170) );
  ND2S U26768 ( .I1(n25258), .I2(n25170), .O(n25171) );
  MUX2 U26769 ( .A(n25171), .B(img[1062]), .S(n29185), .O(n12474) );
  AOI22S U26770 ( .A1(n13781), .A2(n30435), .B1(n28069), .B2(img[1062]), .O(
        n25173) );
  ND3S U26771 ( .I1(n25327), .I2(n25173), .I3(n25172), .O(n25174) );
  MUX2 U26772 ( .A(img[1118]), .B(n25174), .S(n29189), .O(n12414) );
  AOI22S U26773 ( .A1(n29194), .A2(n30436), .B1(n24313), .B2(img[1054]), .O(
        n25176) );
  ND3S U26774 ( .I1(n25327), .I2(n25176), .I3(n25175), .O(n25177) );
  MUX2 U26775 ( .A(img[1126]), .B(n25177), .S(n29198), .O(n12410) );
  AOI22S U26776 ( .A1(n28347), .A2(img[1126]), .B1(n25062), .B2(n30437), .O(
        n25178) );
  ND2S U26777 ( .I1(n25327), .I2(n25178), .O(n25179) );
  AOI22S U26778 ( .A1(n29072), .A2(img[590]), .B1(n28343), .B2(n30438), .O(
        n25180) );
  ND2S U26779 ( .I1(n25327), .I2(n25180), .O(n25181) );
  MUX2 U26780 ( .A(n25181), .B(img[566]), .S(n28578), .O(n12970) );
  AOI22S U26781 ( .A1(n29072), .A2(img[566]), .B1(n13781), .B2(n30439), .O(
        n25182) );
  ND2S U26782 ( .I1(n25327), .I2(n25182), .O(n25183) );
  MUX2 U26783 ( .A(n25183), .B(img[590]), .S(n28581), .O(n12942) );
  AOI22S U26784 ( .A1(n28442), .A2(img[78]), .B1(n13781), .B2(n30440), .O(
        n25184) );
  ND2S U26785 ( .I1(n25327), .I2(n25184), .O(n25185) );
  AOI22S U26786 ( .A1(n28347), .A2(img[54]), .B1(n29407), .B2(n30441), .O(
        n25186) );
  ND2S U26787 ( .I1(n25258), .I2(n25186), .O(n25187) );
  MUX2 U26788 ( .A(img[78]), .B(n25187), .S(n28587), .O(n13454) );
  AOI22S U26789 ( .A1(n25810), .A2(img[974]), .B1(n28135), .B2(n30442), .O(
        n25188) );
  ND2S U26790 ( .I1(n25327), .I2(n25188), .O(n25189) );
  MUX2 U26791 ( .A(n25189), .B(img[950]), .S(n28620), .O(n12582) );
  AOI22S U26792 ( .A1(n28347), .A2(img[950]), .B1(n25591), .B2(n30443), .O(
        n25190) );
  ND2S U26793 ( .I1(n25327), .I2(n25190), .O(n25191) );
  AOI22S U26794 ( .A1(n28106), .A2(img[206]), .B1(n27735), .B2(n30444), .O(
        n25192) );
  ND2S U26795 ( .I1(n25258), .I2(n25192), .O(n25193) );
  MUX2 U26796 ( .A(img[182]), .B(n25193), .S(n28626), .O(n13350) );
  AOI22S U26797 ( .A1(n26970), .A2(img[182]), .B1(n25591), .B2(n30445), .O(
        n25194) );
  ND2S U26798 ( .I1(n25258), .I2(n25194), .O(n25195) );
  MUX2 U26799 ( .A(img[206]), .B(n25195), .S(n28629), .O(n13330) );
  AOI22S U26800 ( .A1(n29072), .A2(img[334]), .B1(n29096), .B2(n30446), .O(
        n25196) );
  ND2S U26801 ( .I1(n25327), .I2(n25196), .O(n25197) );
  MUX2 U26802 ( .A(img[310]), .B(n25197), .S(n28632), .O(n13226) );
  AOI22S U26803 ( .A1(n29435), .A2(img[310]), .B1(n28592), .B2(n30447), .O(
        n25198) );
  ND2S U26804 ( .I1(n25327), .I2(n25198), .O(n25199) );
  AOI22S U26805 ( .A1(n28106), .A2(img[462]), .B1(n13781), .B2(n30448), .O(
        n25200) );
  ND2S U26806 ( .I1(n25258), .I2(n25200), .O(n25201) );
  AOI22S U26807 ( .A1(n24415), .A2(img[438]), .B1(n29242), .B2(n30449), .O(
        n25202) );
  ND2S U26808 ( .I1(n25258), .I2(n25202), .O(n25203) );
  MUX2 U26809 ( .A(n25203), .B(img[462]), .S(n28641), .O(n13074) );
  AOI22S U26810 ( .A1(n28106), .A2(img[846]), .B1(n28433), .B2(n30450), .O(
        n25204) );
  ND2S U26811 ( .I1(n25327), .I2(n25204), .O(n25205) );
  INV1S U26812 ( .I(img[846]), .O(n25206) );
  AOI22S U26813 ( .A1(n29435), .A2(img[822]), .B1(n25591), .B2(n25206), .O(
        n25207) );
  ND2S U26814 ( .I1(n25327), .I2(n25207), .O(n25208) );
  AOI22S U26815 ( .A1(n13771), .A2(img[718]), .B1(n29242), .B2(n30451), .O(
        n25209) );
  ND2S U26816 ( .I1(n25258), .I2(n25209), .O(n25210) );
  AOI22S U26817 ( .A1(n28840), .A2(img[694]), .B1(n25591), .B2(n30452), .O(
        n25211) );
  ND2S U26818 ( .I1(n25327), .I2(n25211), .O(n25212) );
  AOI22S U26819 ( .A1(n29414), .A2(img[606]), .B1(n29096), .B2(n30453), .O(
        n25213) );
  ND2S U26820 ( .I1(n25258), .I2(n25213), .O(n25214) );
  AOI22S U26821 ( .A1(n13778), .A2(img[550]), .B1(n29096), .B2(n30454), .O(
        n25215) );
  ND2S U26822 ( .I1(n25327), .I2(n25215), .O(n25216) );
  MUX2 U26823 ( .A(n25216), .B(img[606]), .S(n29478), .O(n12926) );
  AOI22S U26824 ( .A1(n28840), .A2(img[94]), .B1(n28135), .B2(n30455), .O(
        n25217) );
  ND2S U26825 ( .I1(n25258), .I2(n25217), .O(n25218) );
  MUX2 U26826 ( .A(img[38]), .B(n25218), .S(n29342), .O(n13498) );
  AOI22S U26827 ( .A1(n29072), .A2(img[38]), .B1(n28433), .B2(n30456), .O(
        n25219) );
  ND2S U26828 ( .I1(n25327), .I2(n25219), .O(n25220) );
  AOI22S U26829 ( .A1(n25595), .A2(img[990]), .B1(n25377), .B2(n30457), .O(
        n25221) );
  ND2S U26830 ( .I1(n25327), .I2(n25221), .O(n25222) );
  AOI22S U26831 ( .A1(n28083), .A2(img[934]), .B1(n13781), .B2(n30458), .O(
        n25223) );
  ND2S U26832 ( .I1(n25258), .I2(n25223), .O(n25224) );
  MUX2 U26833 ( .A(img[990]), .B(n25224), .S(n29345), .O(n12546) );
  AOI22S U26834 ( .A1(n13772), .A2(img[222]), .B1(n27511), .B2(n30459), .O(
        n25225) );
  ND2S U26835 ( .I1(n25258), .I2(n25225), .O(n25226) );
  MUX2 U26836 ( .A(img[166]), .B(n25226), .S(n29355), .O(n13366) );
  AOI22S U26837 ( .A1(n28106), .A2(img[166]), .B1(n28075), .B2(n30460), .O(
        n25227) );
  ND2S U26838 ( .I1(n25258), .I2(n25227), .O(n25228) );
  MUX2 U26839 ( .A(img[222]), .B(n25228), .S(n29351), .O(n13314) );
  AOI22S U26840 ( .A1(n25595), .A2(img[350]), .B1(n29407), .B2(n30461), .O(
        n25229) );
  ND2S U26841 ( .I1(n25258), .I2(n25229), .O(n25230) );
  AOI22S U26842 ( .A1(n28442), .A2(img[294]), .B1(n13781), .B2(n30462), .O(
        n25231) );
  ND2S U26843 ( .I1(n25258), .I2(n25231), .O(n25232) );
  MUX2 U26844 ( .A(img[350]), .B(n25232), .S(n29358), .O(n13182) );
  AOI22S U26845 ( .A1(n13776), .A2(img[478]), .B1(n25591), .B2(n30463), .O(
        n25233) );
  ND2S U26846 ( .I1(n25258), .I2(n25233), .O(n25234) );
  MUX2 U26847 ( .A(img[422]), .B(n25234), .S(n29367), .O(n13110) );
  AOI22S U26848 ( .A1(n13773), .A2(img[422]), .B1(n28938), .B2(n30464), .O(
        n25235) );
  ND2S U26849 ( .I1(n25258), .I2(n25235), .O(n25236) );
  MUX2 U26850 ( .A(img[478]), .B(n25236), .S(n29364), .O(n13058) );
  AOI22S U26851 ( .A1(n28347), .A2(img[862]), .B1(n13781), .B2(n30465), .O(
        n25237) );
  ND2S U26852 ( .I1(n25258), .I2(n25237), .O(n25238) );
  MUX2 U26853 ( .A(n25238), .B(img[806]), .S(n29374), .O(n12730) );
  INV1S U26854 ( .I(img[862]), .O(n25239) );
  AOI22S U26855 ( .A1(n28347), .A2(img[806]), .B1(n29242), .B2(n25239), .O(
        n25240) );
  ND2S U26856 ( .I1(n25258), .I2(n25240), .O(n25241) );
  AOI22S U26857 ( .A1(n28840), .A2(img[734]), .B1(n25062), .B2(n30466), .O(
        n25242) );
  ND2S U26858 ( .I1(n25258), .I2(n25242), .O(n25243) );
  AOI22S U26859 ( .A1(n13776), .A2(img[678]), .B1(n28592), .B2(n30467), .O(
        n25244) );
  ND2S U26860 ( .I1(n25258), .I2(n25244), .O(n25245) );
  MUX2 U26861 ( .A(n25245), .B(img[734]), .S(n29377), .O(n12802) );
  AOI22S U26862 ( .A1(n13777), .A2(img[510]), .B1(n24374), .B2(n30468), .O(
        n25246) );
  ND2S U26863 ( .I1(n25258), .I2(n25246), .O(n25247) );
  MUX2 U26864 ( .A(n25247), .B(img[390]), .S(n29416), .O(n13142) );
  INV1S U26865 ( .I(img[510]), .O(n25248) );
  AOI22S U26866 ( .A1(n27990), .A2(img[390]), .B1(n27049), .B2(n25248), .O(
        n25249) );
  ND2S U26867 ( .I1(n25258), .I2(n25249), .O(n25250) );
  AOI22S U26868 ( .A1(n28347), .A2(img[382]), .B1(n13779), .B2(n30469), .O(
        n25251) );
  ND2S U26869 ( .I1(n25258), .I2(n25251), .O(n25252) );
  AOI22S U26870 ( .A1(n13778), .A2(img[262]), .B1(n28433), .B2(n30470), .O(
        n25253) );
  ND2S U26871 ( .I1(n25258), .I2(n25253), .O(n25254) );
  MUX2 U26872 ( .A(img[382]), .B(n25254), .S(n29412), .O(n13150) );
  AOI22S U26873 ( .A1(n27110), .A2(img[638]), .B1(n28695), .B2(n30471), .O(
        n25255) );
  ND2S U26874 ( .I1(n25258), .I2(n25255), .O(n25256) );
  AOI22S U26875 ( .A1(n28840), .A2(img[518]), .B1(n28695), .B2(n30472), .O(
        n25257) );
  ND2S U26876 ( .I1(n25258), .I2(n25257), .O(n25259) );
  MUX2 U26877 ( .A(n25259), .B(img[638]), .S(n29386), .O(n12894) );
  BUF2 U26878 ( .I(n25298), .O(n25338) );
  AOI22S U26879 ( .A1(n27110), .A2(img[126]), .B1(n28433), .B2(n30473), .O(
        n25260) );
  ND2S U26880 ( .I1(n25338), .I2(n25260), .O(n25261) );
  AOI22S U26881 ( .A1(n27110), .A2(img[6]), .B1(n25062), .B2(n30474), .O(
        n25262) );
  ND2S U26882 ( .I1(n25338), .I2(n25262), .O(n25263) );
  MUX2 U26883 ( .A(img[126]), .B(n25263), .S(n29392), .O(n13406) );
  AOI22S U26884 ( .A1(n29072), .A2(img[1022]), .B1(n29530), .B2(n30475), .O(
        n25264) );
  ND2S U26885 ( .I1(n25338), .I2(n25264), .O(n25265) );
  MUX2 U26886 ( .A(img[902]), .B(n25265), .S(n29395), .O(n12630) );
  AOI22S U26887 ( .A1(n26855), .A2(img[902]), .B1(n28433), .B2(n30476), .O(
        n25266) );
  ND2S U26888 ( .I1(n25338), .I2(n25266), .O(n25267) );
  AOI22S U26889 ( .A1(n28347), .A2(img[254]), .B1(n25859), .B2(n30477), .O(
        n25268) );
  ND2S U26890 ( .I1(n25338), .I2(n25268), .O(n25269) );
  MUX2 U26891 ( .A(n25269), .B(img[134]), .S(n29402), .O(n13398) );
  AOI22S U26892 ( .A1(n27990), .A2(img[134]), .B1(n24193), .B2(n30478), .O(
        n25270) );
  ND2S U26893 ( .I1(n25338), .I2(n25270), .O(n25271) );
  MUX2 U26894 ( .A(img[254]), .B(n25271), .S(n29405), .O(n13281) );
  AOI22S U26895 ( .A1(n28347), .A2(img[894]), .B1(n25859), .B2(n30479), .O(
        n25272) );
  ND2S U26896 ( .I1(n25338), .I2(n25272), .O(n25273) );
  MUX2 U26897 ( .A(img[774]), .B(n25273), .S(n29423), .O(n12762) );
  INV1S U26898 ( .I(img[894]), .O(n25274) );
  AOI22S U26899 ( .A1(n29435), .A2(img[774]), .B1(n24193), .B2(n25274), .O(
        n25275) );
  ND2S U26900 ( .I1(n25338), .I2(n25275), .O(n25276) );
  AOI22S U26901 ( .A1(n13777), .A2(img[766]), .B1(n28343), .B2(n30480), .O(
        n25277) );
  ND2S U26902 ( .I1(n25338), .I2(n25277), .O(n25278) );
  AOI22S U26903 ( .A1(n26822), .A2(img[646]), .B1(n25859), .B2(n30481), .O(
        n25279) );
  ND2S U26904 ( .I1(n25338), .I2(n25279), .O(n25280) );
  MUX2 U26905 ( .A(n25280), .B(img[766]), .S(n29433), .O(n12770) );
  AOI22S U26906 ( .A1(n26822), .A2(img[1390]), .B1(n27049), .B2(n30482), .O(
        n25281) );
  ND2S U26907 ( .I1(n25338), .I2(n25281), .O(n25282) );
  MUX2 U26908 ( .A(n25282), .B(img[1302]), .S(n29054), .O(n12234) );
  AOI22S U26909 ( .A1(n25062), .A2(n30483), .B1(n25444), .B2(img[1302]), .O(
        n25284) );
  ND3S U26910 ( .I1(n25327), .I2(n25284), .I3(n25283), .O(n25285) );
  MUX2 U26911 ( .A(img[1390]), .B(n25285), .S(n29058), .O(n12142) );
  AOI22S U26912 ( .A1(n13779), .A2(n30484), .B1(n25444), .B2(img[1326]), .O(
        n25287) );
  ND3S U26913 ( .I1(n25327), .I2(n25287), .I3(n25286), .O(n25288) );
  MUX2 U26914 ( .A(img[1366]), .B(n25288), .S(n29051), .O(n12170) );
  AOI22S U26915 ( .A1(n26822), .A2(img[1366]), .B1(n28343), .B2(n30485), .O(
        n25289) );
  ND2S U26916 ( .I1(n25338), .I2(n25289), .O(n25290) );
  MUX2 U26917 ( .A(n25290), .B(img[1326]), .S(n29047), .O(n12206) );
  AOI22S U26918 ( .A1(n26822), .A2(img[1518]), .B1(n23941), .B2(n30486), .O(
        n25291) );
  ND2S U26919 ( .I1(n25338), .I2(n25291), .O(n25292) );
  AOI22S U26920 ( .A1(n13781), .A2(n30487), .B1(n25444), .B2(img[1430]), .O(
        n25294) );
  ND3S U26921 ( .I1(n25327), .I2(n25294), .I3(n25293), .O(n25295) );
  MUX2 U26922 ( .A(img[1518]), .B(n25295), .S(n29099), .O(n12018) );
  AOI22S U26923 ( .A1(n13781), .A2(n30488), .B1(n25444), .B2(img[1454]), .O(
        n25297) );
  AOI22S U26924 ( .A1(n27110), .A2(img[1494]), .B1(n25062), .B2(n30489), .O(
        n25300) );
  ND2S U26925 ( .I1(n25338), .I2(n25300), .O(n25301) );
  MUX2 U26926 ( .A(n25301), .B(img[1454]), .S(n29087), .O(n12082) );
  AOI22S U26927 ( .A1(n27110), .A2(img[1134]), .B1(n28343), .B2(n30490), .O(
        n25302) );
  ND2S U26928 ( .I1(n25338), .I2(n25302), .O(n25303) );
  MUX2 U26929 ( .A(n25303), .B(img[1046]), .S(n29122), .O(n12489) );
  AOI22S U26930 ( .A1(n28862), .A2(n30491), .B1(n25444), .B2(img[1046]), .O(
        n25305) );
  ND3S U26931 ( .I1(n25327), .I2(n25305), .I3(n25304), .O(n25306) );
  MUX2 U26932 ( .A(img[1134]), .B(n25306), .S(n29127), .O(n12398) );
  AOI22S U26933 ( .A1(n28695), .A2(n30492), .B1(n25444), .B2(img[1070]), .O(
        n25308) );
  ND3S U26934 ( .I1(n25327), .I2(n25308), .I3(n25307), .O(n25309) );
  MUX2 U26935 ( .A(img[1110]), .B(n25309), .S(n29119), .O(n12426) );
  AOI22S U26936 ( .A1(n28840), .A2(img[1110]), .B1(n28433), .B2(n30493), .O(
        n25310) );
  ND2S U26937 ( .I1(n25338), .I2(n25310), .O(n25311) );
  MUX2 U26938 ( .A(n25311), .B(img[1070]), .S(n29115), .O(n12462) );
  AOI22S U26939 ( .A1(n28106), .A2(img[558]), .B1(n25859), .B2(n30494), .O(
        n25312) );
  ND2S U26940 ( .I1(n25338), .I2(n25312), .O(n25313) );
  MUX2 U26941 ( .A(n25313), .B(img[598]), .S(n29133), .O(n12938) );
  AOI22S U26942 ( .A1(n27110), .A2(img[598]), .B1(n25062), .B2(n30495), .O(
        n25314) );
  ND2S U26943 ( .I1(n25338), .I2(n25314), .O(n25315) );
  MUX2 U26944 ( .A(n25315), .B(img[558]), .S(n29439), .O(n12974) );
  AOI22S U26945 ( .A1(n28347), .A2(img[46]), .B1(n28075), .B2(n30496), .O(
        n25316) );
  ND2S U26946 ( .I1(n25338), .I2(n25316), .O(n25317) );
  AOI22S U26947 ( .A1(n27110), .A2(img[86]), .B1(n25062), .B2(n30497), .O(
        n25318) );
  ND2S U26948 ( .I1(n25338), .I2(n25318), .O(n25319) );
  MUX2 U26949 ( .A(img[46]), .B(n25319), .S(n29136), .O(n13486) );
  AOI22S U26950 ( .A1(n26855), .A2(img[1262]), .B1(n25859), .B2(n30498), .O(
        n25320) );
  ND2S U26951 ( .I1(n25338), .I2(n25320), .O(n25321) );
  AOI22S U26952 ( .A1(n28343), .A2(n30499), .B1(n25444), .B2(img[1174]), .O(
        n25323) );
  ND3S U26953 ( .I1(n25327), .I2(n25323), .I3(n25322), .O(n25324) );
  MUX2 U26954 ( .A(img[1262]), .B(n25324), .S(n29044), .O(n12274) );
  AOI22S U26955 ( .A1(n28135), .A2(n30500), .B1(n25444), .B2(img[1198]), .O(
        n25326) );
  ND3S U26956 ( .I1(n25327), .I2(n25326), .I3(n25325), .O(n25328) );
  MUX2 U26957 ( .A(img[1238]), .B(n25328), .S(n29037), .O(n12294) );
  AOI22S U26958 ( .A1(n26855), .A2(img[1238]), .B1(n25859), .B2(n30501), .O(
        n25329) );
  ND2S U26959 ( .I1(n25338), .I2(n25329), .O(n25330) );
  MUX2 U26960 ( .A(img[1198]), .B(n25330), .S(n29033), .O(n12338) );
  AOI22S U26961 ( .A1(n25810), .A2(img[942]), .B1(n25062), .B2(n30502), .O(
        n25331) );
  ND2S U26962 ( .I1(n25338), .I2(n25331), .O(n25332) );
  MUX2 U26963 ( .A(img[982]), .B(n25332), .S(n29145), .O(n12550) );
  AOI22S U26964 ( .A1(n28347), .A2(img[982]), .B1(n24193), .B2(n30503), .O(
        n25333) );
  ND2S U26965 ( .I1(n25338), .I2(n25333), .O(n25334) );
  AOI22S U26966 ( .A1(n26822), .A2(img[174]), .B1(n28695), .B2(n30504), .O(
        n25335) );
  ND2S U26967 ( .I1(n25338), .I2(n25335), .O(n25336) );
  MUX2 U26968 ( .A(img[214]), .B(n25336), .S(n29151), .O(n13318) );
  AOI22S U26969 ( .A1(n26822), .A2(img[214]), .B1(n28695), .B2(n30505), .O(
        n25337) );
  ND2S U26970 ( .I1(n25338), .I2(n25337), .O(n25339) );
  MUX2 U26971 ( .A(img[174]), .B(n25339), .S(n29148), .O(n13362) );
  AOI22S U26972 ( .A1(n26822), .A2(img[302]), .B1(n25062), .B2(n30506), .O(
        n25340) );
  ND2S U26973 ( .I1(n25327), .I2(n25340), .O(n25341) );
  MUX2 U26974 ( .A(img[342]), .B(n25341), .S(n29157), .O(n13194) );
  AOI22S U26975 ( .A1(n26822), .A2(img[342]), .B1(n24193), .B2(n30507), .O(
        n25342) );
  ND2S U26976 ( .I1(n25327), .I2(n25342), .O(n25343) );
  AOI22S U26977 ( .A1(n26822), .A2(img[430]), .B1(n25062), .B2(n30508), .O(
        n25344) );
  ND2S U26978 ( .I1(n25327), .I2(n25344), .O(n25345) );
  MUX2 U26979 ( .A(img[470]), .B(n25345), .S(n29163), .O(n13062) );
  AOI22S U26980 ( .A1(n26822), .A2(img[470]), .B1(n23918), .B2(n30509), .O(
        n25346) );
  ND2S U26981 ( .I1(n25327), .I2(n25346), .O(n25347) );
  MUX2 U26982 ( .A(img[430]), .B(n25347), .S(n29160), .O(n13106) );
  INV1S U26983 ( .I(img[854]), .O(n25348) );
  AOI22S U26984 ( .A1(n26822), .A2(img[814]), .B1(n28037), .B2(n25348), .O(
        n25349) );
  ND2S U26985 ( .I1(n25327), .I2(n25349), .O(n25350) );
  AOI22S U26986 ( .A1(n13772), .A2(img[854]), .B1(n13781), .B2(n30510), .O(
        n25351) );
  ND2S U26987 ( .I1(n25327), .I2(n25351), .O(n25352) );
  MUX2 U26988 ( .A(n25352), .B(img[814]), .S(n29166), .O(n12718) );
  AOI22S U26989 ( .A1(n29072), .A2(img[686]), .B1(n25591), .B2(n30511), .O(
        n25353) );
  ND2S U26990 ( .I1(n25327), .I2(n25353), .O(n25354) );
  AOI22S U26991 ( .A1(n13778), .A2(img[726]), .B1(n25062), .B2(n30512), .O(
        n25355) );
  ND2S U26992 ( .I1(n25327), .I2(n25355), .O(n25356) );
  AOI22S U26993 ( .A1(n29414), .A2(img[622]), .B1(n24755), .B2(n30513), .O(
        n25357) );
  ND2S U26994 ( .I1(n25327), .I2(n25357), .O(n25358) );
  AOI22S U26995 ( .A1(n29435), .A2(img[534]), .B1(n25591), .B2(n30514), .O(
        n25359) );
  ND2S U26996 ( .I1(n25327), .I2(n25359), .O(n25360) );
  MUX2 U26997 ( .A(n25360), .B(img[622]), .S(n29024), .O(n12910) );
  AOI22S U26998 ( .A1(n13773), .A2(img[110]), .B1(n25062), .B2(n30515), .O(
        n25361) );
  ND2S U26999 ( .I1(n25327), .I2(n25361), .O(n25362) );
  MUX2 U27000 ( .A(img[22]), .B(n25362), .S(n29027), .O(n13514) );
  AOI22S U27001 ( .A1(n26970), .A2(img[22]), .B1(n29096), .B2(n30516), .O(
        n25363) );
  ND2S U27002 ( .I1(n25327), .I2(n25363), .O(n25364) );
  AOI22S U27003 ( .A1(n28318), .A2(img[1006]), .B1(n29096), .B2(n30517), .O(
        n25365) );
  ND2S U27004 ( .I1(n25327), .I2(n25365), .O(n25366) );
  MUX2 U27005 ( .A(img[918]), .B(n25366), .S(n29061), .O(n12614) );
  AOI22S U27006 ( .A1(n27990), .A2(img[918]), .B1(n28614), .B2(n30518), .O(
        n25367) );
  ND2S U27007 ( .I1(n25327), .I2(n25367), .O(n25368) );
  AOI22S U27008 ( .A1(n28347), .A2(img[238]), .B1(n13775), .B2(n30519), .O(
        n25369) );
  ND2S U27009 ( .I1(n25327), .I2(n25369), .O(n25370) );
  AOI22S U27010 ( .A1(n28382), .A2(img[150]), .B1(n25062), .B2(n30520), .O(
        n25371) );
  ND2S U27011 ( .I1(n25327), .I2(n25371), .O(n25372) );
  MUX2 U27012 ( .A(img[238]), .B(n25372), .S(n29070), .O(n13298) );
  AOI22S U27013 ( .A1(n28318), .A2(img[366]), .B1(n28614), .B2(n30521), .O(
        n25373) );
  ND2S U27014 ( .I1(n25327), .I2(n25373), .O(n25374) );
  AOI22S U27015 ( .A1(n28347), .A2(img[278]), .B1(n28695), .B2(n30522), .O(
        n25375) );
  ND2S U27016 ( .I1(n25327), .I2(n25375), .O(n25376) );
  MUX2 U27017 ( .A(img[366]), .B(n25376), .S(n29078), .O(n13166) );
  AOI22S U27018 ( .A1(n26855), .A2(img[494]), .B1(n27049), .B2(n30523), .O(
        n25378) );
  ND2S U27019 ( .I1(n25327), .I2(n25378), .O(n25379) );
  AOI22S U27020 ( .A1(n28347), .A2(img[406]), .B1(n28037), .B2(n30524), .O(
        n25380) );
  ND2S U27021 ( .I1(n25327), .I2(n25380), .O(n25381) );
  MUX2 U27022 ( .A(img[494]), .B(n25381), .S(n29084), .O(n13042) );
  AOI22S U27023 ( .A1(n29414), .A2(img[878]), .B1(n28162), .B2(n30525), .O(
        n25382) );
  ND2S U27024 ( .I1(n25327), .I2(n25382), .O(n25383) );
  MUX2 U27025 ( .A(img[790]), .B(n25383), .S(n29102), .O(n12746) );
  INV1S U27026 ( .I(img[878]), .O(n25384) );
  AOI22S U27027 ( .A1(n13772), .A2(img[790]), .B1(n28075), .B2(n25384), .O(
        n25385) );
  ND2S U27028 ( .I1(n25327), .I2(n25385), .O(n25386) );
  AOI22S U27029 ( .A1(n26855), .A2(img[750]), .B1(n29530), .B2(n30526), .O(
        n25387) );
  ND2S U27030 ( .I1(n25327), .I2(n25387), .O(n25388) );
  AOI22S U27031 ( .A1(n28442), .A2(img[662]), .B1(n29194), .B2(n30527), .O(
        n25389) );
  ND2S U27032 ( .I1(n25327), .I2(n25389), .O(n25390) );
  OAI22S U27033 ( .A1(n25392), .A2(n28530), .B1(n13897), .B2(n25391), .O(
        n25393) );
  AOI12HS U27034 ( .B1(n28534), .B2(n29484), .A1(n25393), .O(n25394) );
  ND2S U27035 ( .I1(n28547), .I2(A67_shift[250]), .O(n25398) );
  AOI22S U27036 ( .A1(n28550), .A2(A67_shift[90]), .B1(n28551), .B2(
        A67_shift[218]), .O(n25397) );
  ND2S U27037 ( .I1(n28554), .I2(A67_shift[122]), .O(n25396) );
  INV1S U27038 ( .I(A67_shift[58]), .O(n25401) );
  AOI22S U27039 ( .A1(n28553), .A2(A67_shift[26]), .B1(n28546), .B2(
        A67_shift[186]), .O(n25400) );
  AOI12HS U27040 ( .B1(n28552), .B2(A67_shift[154]), .A1(n28555), .O(n25399)
         );
  OAI112HS U27041 ( .C1(n28544), .C2(n25401), .A1(n25400), .B1(n25399), .O(
        n25413) );
  INV1S U27042 ( .I(A67_shift[42]), .O(n25402) );
  NR2 U27043 ( .I1(n25402), .I2(n28544), .O(n25408) );
  ND2S U27044 ( .I1(n28552), .I2(A67_shift[138]), .O(n25404) );
  ND2S U27045 ( .I1(A67_shift[234]), .I2(n28547), .O(n25403) );
  INV1S U27046 ( .I(A67_shift[170]), .O(n25405) );
  MOAI1S U27047 ( .A1(n26653), .A2(n25405), .B1(n28551), .B2(A67_shift[202]), 
        .O(n25406) );
  NR3 U27048 ( .I1(n25408), .I2(n25407), .I3(n25406), .O(n25411) );
  AOI22S U27049 ( .A1(n28550), .A2(A67_shift[74]), .B1(n28553), .B2(
        A67_shift[10]), .O(n25410) );
  OAI12HS U27050 ( .B1(n25414), .B2(n25413), .A1(n25412), .O(n25418) );
  AOI22S U27051 ( .A1(n28566), .A2(gray_max_out[2]), .B1(n28565), .B2(
        gray_weight_out[2]), .O(n25416) );
  ND2S U27052 ( .I1(n28564), .I2(gray_avg_out[2]), .O(n25415) );
  AOI22S U27053 ( .A1(n28382), .A2(img[522]), .B1(n28343), .B2(n30528), .O(
        n25421) );
  ND2S U27054 ( .I1(n26010), .I2(n25421), .O(n25422) );
  MUX2 U27055 ( .A(n25422), .B(img[626]), .S(n29292), .O(n12902) );
  AOI22S U27056 ( .A1(n27746), .A2(img[626]), .B1(n28135), .B2(n30529), .O(
        n25423) );
  ND2S U27057 ( .I1(n26010), .I2(n25423), .O(n25424) );
  AOI22S U27058 ( .A1(n28382), .A2(img[10]), .B1(n25591), .B2(n30530), .O(
        n25425) );
  ND2S U27059 ( .I1(n26010), .I2(n25425), .O(n25426) );
  AOI22S U27060 ( .A1(n13773), .A2(img[114]), .B1(n27049), .B2(n30531), .O(
        n25427) );
  ND2S U27061 ( .I1(n26010), .I2(n25427), .O(n25428) );
  MUX2 U27062 ( .A(n25428), .B(img[10]), .S(n29295), .O(n13522) );
  AOI22S U27063 ( .A1(n13773), .A2(img[1226]), .B1(n27511), .B2(n30532), .O(
        n25429) );
  ND2S U27064 ( .I1(n26010), .I2(n25429), .O(n25430) );
  AOI22S U27065 ( .A1(n28938), .A2(n30533), .B1(n25444), .B2(img[1202]), .O(
        n25432) );
  ND3S U27066 ( .I1(n26010), .I2(n25432), .I3(n25431), .O(n25433) );
  MUX2 U27067 ( .A(img[1226]), .B(n25433), .S(n28602), .O(n12302) );
  AOI22S U27068 ( .A1(n28075), .A2(n30534), .B1(n25444), .B2(img[1162]), .O(
        n25435) );
  ND3S U27069 ( .I1(n26010), .I2(n25435), .I3(n25434), .O(n25436) );
  MUX2 U27070 ( .A(img[1266]), .B(n25436), .S(n28595), .O(n12266) );
  AOI22S U27071 ( .A1(n13773), .A2(img[1266]), .B1(n28433), .B2(n30535), .O(
        n25437) );
  ND2S U27072 ( .I1(n26010), .I2(n25437), .O(n25438) );
  AOI22S U27073 ( .A1(n13773), .A2(img[1354]), .B1(n29242), .B2(n30536), .O(
        n25439) );
  ND2S U27074 ( .I1(n26010), .I2(n25439), .O(n25440) );
  MUX2 U27075 ( .A(n25440), .B(img[1330]), .S(n28612), .O(n12198) );
  AOI22S U27076 ( .A1(n28592), .A2(n30537), .B1(n25444), .B2(img[1330]), .O(
        n25442) );
  ND3S U27077 ( .I1(n26010), .I2(n25442), .I3(n25441), .O(n25443) );
  MUX2 U27078 ( .A(img[1354]), .B(n25443), .S(n28617), .O(n12178) );
  AOI22S U27079 ( .A1(n28162), .A2(n30538), .B1(n25444), .B2(img[1290]), .O(
        n25446) );
  ND3S U27080 ( .I1(n26010), .I2(n25446), .I3(n25445), .O(n25447) );
  MUX2 U27081 ( .A(img[1394]), .B(n25447), .S(n28609), .O(n12134) );
  AOI22S U27082 ( .A1(n28382), .A2(img[1394]), .B1(n29242), .B2(n30539), .O(
        n25448) );
  ND2S U27083 ( .I1(n26010), .I2(n25448), .O(n25449) );
  AOI22S U27084 ( .A1(n13776), .A2(img[906]), .B1(n29096), .B2(n30540), .O(
        n25450) );
  ND2S U27085 ( .I1(n26010), .I2(n25450), .O(n25451) );
  AOI22S U27086 ( .A1(n28083), .A2(img[1010]), .B1(n25062), .B2(n30541), .O(
        n25452) );
  ND2S U27087 ( .I1(n26010), .I2(n25452), .O(n25453) );
  MUX2 U27088 ( .A(img[906]), .B(n25453), .S(n29300), .O(n12622) );
  AOI22S U27089 ( .A1(n13772), .A2(img[138]), .B1(n27443), .B2(n30542), .O(
        n25454) );
  ND2S U27090 ( .I1(n26010), .I2(n25454), .O(n25455) );
  MUX2 U27091 ( .A(img[242]), .B(n25455), .S(n29309), .O(n13290) );
  AOI22S U27092 ( .A1(n28382), .A2(img[242]), .B1(n28182), .B2(n30543), .O(
        n25456) );
  ND2S U27093 ( .I1(n26010), .I2(n25456), .O(n25457) );
  MUX2 U27094 ( .A(img[138]), .B(n25457), .S(n29306), .O(n13390) );
  AOI22S U27095 ( .A1(n28382), .A2(img[266]), .B1(n28592), .B2(n30544), .O(
        n25458) );
  ND2S U27096 ( .I1(n26010), .I2(n25458), .O(n25459) );
  AOI22S U27097 ( .A1(n28347), .A2(img[370]), .B1(n23918), .B2(n30545), .O(
        n25460) );
  ND2S U27098 ( .I1(n26010), .I2(n25460), .O(n25461) );
  MUX2 U27099 ( .A(n25461), .B(img[266]), .S(n29312), .O(n13266) );
  AOI22S U27100 ( .A1(n13776), .A2(img[394]), .B1(n29457), .B2(n30546), .O(
        n25462) );
  ND2S U27101 ( .I1(n26010), .I2(n25462), .O(n25463) );
  AOI22S U27102 ( .A1(n13776), .A2(img[498]), .B1(n29397), .B2(n30547), .O(
        n25464) );
  ND2S U27103 ( .I1(n26010), .I2(n25464), .O(n25465) );
  MUX2 U27104 ( .A(n25465), .B(img[394]), .S(n29318), .O(n13134) );
  AOI22S U27105 ( .A1(n13776), .A2(img[1482]), .B1(n13779), .B2(n30548), .O(
        n25466) );
  ND2S U27106 ( .I1(n26010), .I2(n25466), .O(n25467) );
  MUX2 U27107 ( .A(img[1458]), .B(n25467), .S(n28652), .O(n12074) );
  BUF12CK U27108 ( .I(n25903), .O(n26010) );
  AOI22S U27109 ( .A1(n25591), .A2(n30549), .B1(n24434), .B2(img[1458]), .O(
        n25470) );
  ND3S U27110 ( .I1(n26010), .I2(n25470), .I3(n25469), .O(n25471) );
  MUX2 U27111 ( .A(img[1482]), .B(n25471), .S(n28656), .O(n12046) );
  AOI22S U27112 ( .A1(n29407), .A2(n30550), .B1(n24946), .B2(img[1418]), .O(
        n25473) );
  ND3S U27113 ( .I1(n26010), .I2(n25473), .I3(n25472), .O(n25474) );
  MUX2 U27114 ( .A(img[1522]), .B(n25474), .S(n28649), .O(n12010) );
  AOI22S U27115 ( .A1(n13776), .A2(img[1522]), .B1(n24193), .B2(n30551), .O(
        n25475) );
  ND2S U27116 ( .I1(n26010), .I2(n25475), .O(n25476) );
  INV1S U27117 ( .I(img[882]), .O(n25477) );
  AOI22S U27118 ( .A1(n13773), .A2(img[778]), .B1(n27049), .B2(n25477), .O(
        n25478) );
  ND2S U27119 ( .I1(n26010), .I2(n25478), .O(n25479) );
  AOI22S U27120 ( .A1(n13773), .A2(img[882]), .B1(n27049), .B2(n30552), .O(
        n25480) );
  ND2S U27121 ( .I1(n26010), .I2(n25480), .O(n25481) );
  MUX2 U27122 ( .A(img[778]), .B(n25481), .S(n29324), .O(n12754) );
  AOI22S U27123 ( .A1(n13773), .A2(img[650]), .B1(n29457), .B2(n30553), .O(
        n25482) );
  ND2S U27124 ( .I1(n26010), .I2(n25482), .O(n25483) );
  AOI22S U27125 ( .A1(n13773), .A2(img[754]), .B1(n29407), .B2(n30554), .O(
        n25484) );
  ND2S U27126 ( .I1(n26010), .I2(n25484), .O(n25485) );
  AOI22S U27127 ( .A1(n13773), .A2(img[1874]), .B1(n29457), .B2(n30555), .O(
        n25486) );
  ND2S U27128 ( .I1(n26010), .I2(n25486), .O(n25487) );
  MUX2 U27129 ( .A(n25487), .B(img[1834]), .S(n28672), .O(n11698) );
  AOI22S U27130 ( .A1(n28135), .A2(n30556), .B1(n24313), .B2(img[1834]), .O(
        n25489) );
  ND2S U27131 ( .I1(n13770), .I2(img[1898]), .O(n25488) );
  ND3S U27132 ( .I1(n26010), .I2(n25489), .I3(n25488), .O(n25490) );
  MUX2 U27133 ( .A(img[1874]), .B(n25490), .S(n28676), .O(n11654) );
  AOI22S U27134 ( .A1(n13773), .A2(img[1898]), .B1(n25591), .B2(n30557), .O(
        n25491) );
  ND2S U27135 ( .I1(n26010), .I2(n25491), .O(n25492) );
  MUX2 U27136 ( .A(n25492), .B(img[1810]), .S(n28679), .O(n11718) );
  AOI22S U27137 ( .A1(n28862), .A2(n30558), .B1(n24313), .B2(img[1810]), .O(
        n25494) );
  AOI22S U27138 ( .A1(n29124), .A2(img[1874]), .B1(img[1906]), .B2(n13782), 
        .O(n25493) );
  ND3S U27139 ( .I1(n26010), .I2(n25494), .I3(n25493), .O(n25495) );
  MUX2 U27140 ( .A(img[1898]), .B(n25495), .S(n28683), .O(n11634) );
  AOI22S U27141 ( .A1(n13773), .A2(img[1866]), .B1(n25377), .B2(n30559), .O(
        n25496) );
  ND2S U27142 ( .I1(n26010), .I2(n25496), .O(n25497) );
  MUX2 U27143 ( .A(n25497), .B(img[1842]), .S(n28693), .O(n11686) );
  AOI22S U27144 ( .A1(n28182), .A2(n30560), .B1(n24313), .B2(img[1842]), .O(
        n25499) );
  ND3S U27145 ( .I1(n26010), .I2(n25499), .I3(n25498), .O(n25500) );
  MUX2 U27146 ( .A(img[1866]), .B(n25500), .S(n28698), .O(n11666) );
  AOI22S U27147 ( .A1(n28182), .A2(n30561), .B1(n24946), .B2(img[1802]), .O(
        n25502) );
  AOI22S U27148 ( .A1(n13905), .A2(img[1866]), .B1(img[1898]), .B2(n28908), 
        .O(n25501) );
  ND3S U27149 ( .I1(n26010), .I2(n25502), .I3(n25501), .O(n25503) );
  MUX2 U27150 ( .A(img[1906]), .B(n25503), .S(n28690), .O(n11622) );
  AOI22S U27151 ( .A1(n25595), .A2(img[1906]), .B1(n25377), .B2(n30562), .O(
        n25504) );
  ND2S U27152 ( .I1(n26010), .I2(n25504), .O(n25505) );
  AOI22S U27153 ( .A1(n25595), .A2(img[1746]), .B1(n28862), .B2(n30563), .O(
        n25506) );
  ND2S U27154 ( .I1(n26010), .I2(n25506), .O(n25507) );
  AOI22S U27155 ( .A1(n28037), .A2(n30564), .B1(n28069), .B2(img[1706]), .O(
        n25509) );
  ND2S U27156 ( .I1(n13770), .I2(img[1770]), .O(n25508) );
  ND3S U27157 ( .I1(n26010), .I2(n25509), .I3(n25508), .O(n25510) );
  MUX2 U27158 ( .A(img[1746]), .B(n25510), .S(n28705), .O(n11786) );
  AOI22S U27159 ( .A1(n25595), .A2(img[1770]), .B1(n28913), .B2(n30565), .O(
        n25511) );
  ND2S U27160 ( .I1(n13769), .I2(n25511), .O(n25512) );
  AOI22S U27161 ( .A1(n28037), .A2(n30566), .B1(n28069), .B2(img[1682]), .O(
        n25514) );
  AOI22S U27162 ( .A1(n13903), .A2(img[1746]), .B1(img[1778]), .B2(n28908), 
        .O(n25513) );
  ND3S U27163 ( .I1(n26010), .I2(n25514), .I3(n25513), .O(n25515) );
  MUX2 U27164 ( .A(img[1770]), .B(n25515), .S(n28712), .O(n11758) );
  AOI22S U27165 ( .A1(n25595), .A2(img[1738]), .B1(n27511), .B2(n30567), .O(
        n25516) );
  ND2S U27166 ( .I1(n26010), .I2(n25516), .O(n25517) );
  MUX2 U27167 ( .A(n25517), .B(img[1714]), .S(n28722), .O(n11818) );
  AOI22S U27168 ( .A1(n28037), .A2(n30568), .B1(n29257), .B2(img[1714]), .O(
        n25519) );
  ND2S U27169 ( .I1(n29258), .I2(img[1778]), .O(n25518) );
  ND3S U27170 ( .I1(n26010), .I2(n25519), .I3(n25518), .O(n25520) );
  MUX2 U27171 ( .A(img[1738]), .B(n25520), .S(n28726), .O(n11790) );
  AOI22S U27172 ( .A1(n28162), .A2(n30569), .B1(n24808), .B2(img[1674]), .O(
        n25522) );
  AOI22S U27173 ( .A1(n13900), .A2(img[1738]), .B1(img[1770]), .B2(n13782), 
        .O(n25521) );
  ND3S U27174 ( .I1(n26010), .I2(n25522), .I3(n25521), .O(n25523) );
  MUX2 U27175 ( .A(img[1778]), .B(n25523), .S(n28719), .O(n11754) );
  AOI22S U27176 ( .A1(n13776), .A2(img[1778]), .B1(n27511), .B2(n30570), .O(
        n25524) );
  ND2S U27177 ( .I1(n26010), .I2(n25524), .O(n25525) );
  AOI22S U27178 ( .A1(n13776), .A2(img[1618]), .B1(n27511), .B2(n30571), .O(
        n25526) );
  ND2S U27179 ( .I1(n26010), .I2(n25526), .O(n25527) );
  MUX2 U27180 ( .A(n25527), .B(img[1578]), .S(n28729), .O(n11954) );
  AOI22S U27181 ( .A1(n28162), .A2(n30572), .B1(n24946), .B2(img[1578]), .O(
        n25529) );
  ND2S U27182 ( .I1(n13770), .I2(img[1642]), .O(n25528) );
  ND3S U27183 ( .I1(n26010), .I2(n25529), .I3(n25528), .O(n25530) );
  MUX2 U27184 ( .A(img[1618]), .B(n25530), .S(n28733), .O(n11910) );
  AOI22S U27185 ( .A1(n13776), .A2(img[1642]), .B1(n13775), .B2(n30573), .O(
        n25531) );
  ND2S U27186 ( .I1(n26010), .I2(n25531), .O(n25532) );
  MUX2 U27187 ( .A(n25532), .B(img[1554]), .S(n28736), .O(n11974) );
  AOI22S U27188 ( .A1(n28162), .A2(n30574), .B1(n24808), .B2(img[1554]), .O(
        n25534) );
  AOI22S U27189 ( .A1(n13904), .A2(img[1618]), .B1(img[1650]), .B2(n13782), 
        .O(n25533) );
  ND3S U27190 ( .I1(n26010), .I2(n25534), .I3(n25533), .O(n25535) );
  MUX2 U27191 ( .A(img[1642]), .B(n25535), .S(n28740), .O(n11890) );
  AOI22S U27192 ( .A1(n13776), .A2(img[1610]), .B1(n24374), .B2(n30575), .O(
        n25536) );
  ND2S U27193 ( .I1(n13769), .I2(n25536), .O(n25537) );
  AOI22S U27194 ( .A1(n28182), .A2(n30576), .B1(n28069), .B2(img[1586]), .O(
        n25539) );
  ND2S U27195 ( .I1(n13770), .I2(img[1650]), .O(n25538) );
  ND3S U27196 ( .I1(n26010), .I2(n25539), .I3(n25538), .O(n25540) );
  MUX2 U27197 ( .A(img[1610]), .B(n25540), .S(n28754), .O(n11922) );
  AOI22S U27198 ( .A1(n28162), .A2(n30577), .B1(n28069), .B2(img[1546]), .O(
        n25542) );
  AOI22S U27199 ( .A1(n13770), .A2(img[1610]), .B1(img[1642]), .B2(n13782), 
        .O(n25541) );
  ND3S U27200 ( .I1(n26010), .I2(n25542), .I3(n25541), .O(n25543) );
  MUX2 U27201 ( .A(img[1650]), .B(n25543), .S(n28747), .O(n11878) );
  AOI22S U27202 ( .A1(n13776), .A2(img[1650]), .B1(n28614), .B2(n30578), .O(
        n25544) );
  ND2S U27203 ( .I1(n26010), .I2(n25544), .O(n25545) );
  AOI22S U27204 ( .A1(n13776), .A2(img[1098]), .B1(n28862), .B2(n30579), .O(
        n25546) );
  ND2S U27205 ( .I1(n26010), .I2(n25546), .O(n25547) );
  MUX2 U27206 ( .A(n25547), .B(img[1074]), .S(n28764), .O(n12454) );
  AOI22S U27207 ( .A1(n28162), .A2(n30580), .B1(n28069), .B2(img[1074]), .O(
        n25549) );
  ND3S U27208 ( .I1(n26010), .I2(n25549), .I3(n25548), .O(n25550) );
  MUX2 U27209 ( .A(img[1098]), .B(n25550), .S(n28768), .O(n12434) );
  AOI22S U27210 ( .A1(n25591), .A2(n30581), .B1(n25444), .B2(img[1034]), .O(
        n25552) );
  ND2S U27211 ( .I1(n29124), .I2(img[1098]), .O(n25551) );
  AOI22S U27212 ( .A1(n13776), .A2(img[1138]), .B1(n24755), .B2(n30582), .O(
        n25554) );
  ND2S U27213 ( .I1(n26010), .I2(n25554), .O(n25555) );
  AOI22S U27214 ( .A1(n25810), .A2(img[2002]), .B1(n13779), .B2(n30583), .O(
        n25556) );
  ND2S U27215 ( .I1(n26010), .I2(n25556), .O(n25557) );
  MUX2 U27216 ( .A(n25557), .B(img[1962]), .S(n28771), .O(n11566) );
  AOI22S U27217 ( .A1(n25377), .A2(n30584), .B1(n25444), .B2(img[1962]), .O(
        n25559) );
  ND3S U27218 ( .I1(n26010), .I2(n25559), .I3(n25558), .O(n25560) );
  MUX2 U27219 ( .A(img[2002]), .B(n25560), .S(n28775), .O(n11530) );
  AOI22S U27220 ( .A1(n28468), .A2(img[2026]), .B1(n13779), .B2(n30585), .O(
        n25561) );
  ND2S U27221 ( .I1(n26010), .I2(n25561), .O(n25562) );
  MUX2 U27222 ( .A(n25562), .B(img[1938]), .S(n28778), .O(n11594) );
  AOI22S U27223 ( .A1(n24193), .A2(n30586), .B1(n24313), .B2(img[1938]), .O(
        n25564) );
  AOI22S U27224 ( .A1(n13903), .A2(img[2002]), .B1(img[2034]), .B2(n13782), 
        .O(n25563) );
  ND3 U27225 ( .I1(n25903), .I2(n25564), .I3(n25563), .O(n25565) );
  AOI22S U27226 ( .A1(n13771), .A2(img[1994]), .B1(n13779), .B2(n30587), .O(
        n25566) );
  ND2S U27227 ( .I1(n26010), .I2(n25566), .O(n25567) );
  MUX2 U27228 ( .A(n25567), .B(img[1970]), .S(n28792), .O(n11562) );
  AOI22S U27229 ( .A1(n23941), .A2(n30588), .B1(n28069), .B2(img[1970]), .O(
        n25569) );
  ND3S U27230 ( .I1(n26010), .I2(n25569), .I3(n25568), .O(n25570) );
  MUX2 U27231 ( .A(img[1994]), .B(n25570), .S(n28796), .O(n11534) );
  AOI22S U27232 ( .A1(n27735), .A2(n30589), .B1(n27919), .B2(img[1930]), .O(
        n25572) );
  AOI22S U27233 ( .A1(n13899), .A2(img[1994]), .B1(img[2026]), .B2(n28908), 
        .O(n25571) );
  ND3S U27234 ( .I1(n26010), .I2(n25572), .I3(n25571), .O(n25573) );
  MUX2 U27235 ( .A(img[2034]), .B(n25573), .S(n28789), .O(n11498) );
  AOI22S U27236 ( .A1(n27065), .A2(img[2034]), .B1(n13779), .B2(n30590), .O(
        n25574) );
  ND2S U27237 ( .I1(n26010), .I2(n25574), .O(n25575) );
  MUX2 U27238 ( .A(img[1930]), .B(n25575), .S(n28785), .O(n11598) );
  AOI22S U27239 ( .A1(n25595), .A2(img[594]), .B1(n27511), .B2(n30591), .O(
        n25576) );
  ND2S U27240 ( .I1(n26010), .I2(n25576), .O(n25577) );
  MUX2 U27241 ( .A(n25577), .B(img[554]), .S(n29439), .O(n12978) );
  AOI22S U27242 ( .A1(n25595), .A2(img[554]), .B1(n27049), .B2(n30592), .O(
        n25578) );
  ND2S U27243 ( .I1(n26010), .I2(n25578), .O(n25579) );
  MUX2 U27244 ( .A(n25579), .B(img[594]), .S(n29133), .O(n12934) );
  AOI22S U27245 ( .A1(n25595), .A2(img[82]), .B1(n27049), .B2(n30593), .O(
        n25580) );
  ND2S U27246 ( .I1(n26010), .I2(n25580), .O(n25581) );
  MUX2 U27247 ( .A(img[42]), .B(n25581), .S(n29136), .O(n13490) );
  AOI22S U27248 ( .A1(n25595), .A2(img[42]), .B1(n27049), .B2(n30594), .O(
        n25582) );
  ND2S U27249 ( .I1(n26010), .I2(n25582), .O(n25583) );
  AOI22S U27250 ( .A1(n25595), .A2(img[1258]), .B1(n27049), .B2(n30595), .O(
        n25584) );
  ND2S U27251 ( .I1(n26010), .I2(n25584), .O(n25585) );
  MUX2 U27252 ( .A(img[1170]), .B(n25585), .S(n29040), .O(n12362) );
  AOI22S U27253 ( .A1(n28135), .A2(n30596), .B1(n24946), .B2(img[1170]), .O(
        n25587) );
  ND3S U27254 ( .I1(n26010), .I2(n25587), .I3(n25586), .O(n25588) );
  MUX2 U27255 ( .A(img[1258]), .B(n25588), .S(n29044), .O(n12270) );
  AOI22S U27256 ( .A1(n25595), .A2(img[1234]), .B1(n28182), .B2(n30597), .O(
        n25589) );
  ND2S U27257 ( .I1(n26010), .I2(n25589), .O(n25590) );
  AOI22S U27258 ( .A1(n27735), .A2(n30598), .B1(n28069), .B2(img[1194]), .O(
        n25593) );
  ND2S U27259 ( .I1(n29124), .I2(img[1258]), .O(n25592) );
  ND3S U27260 ( .I1(n26010), .I2(n25593), .I3(n25592), .O(n25594) );
  MUX2 U27261 ( .A(img[1234]), .B(n25594), .S(n29037), .O(n12298) );
  AOI22S U27262 ( .A1(n25595), .A2(img[1386]), .B1(n28182), .B2(n30599), .O(
        n25596) );
  ND2S U27263 ( .I1(n26010), .I2(n25596), .O(n25597) );
  MUX2 U27264 ( .A(n25597), .B(img[1298]), .S(n29054), .O(n12230) );
  AOI22S U27265 ( .A1(n25377), .A2(n30600), .B1(n25444), .B2(img[1298]), .O(
        n25599) );
  ND3S U27266 ( .I1(n26010), .I2(n25599), .I3(n25598), .O(n25600) );
  MUX2 U27267 ( .A(img[1386]), .B(n25600), .S(n29058), .O(n12146) );
  AOI22S U27268 ( .A1(n13777), .A2(img[1362]), .B1(n28162), .B2(n30601), .O(
        n25601) );
  ND2S U27269 ( .I1(n26010), .I2(n25601), .O(n25602) );
  AOI22S U27270 ( .A1(n25377), .A2(n30602), .B1(n24313), .B2(img[1322]), .O(
        n25604) );
  ND2S U27271 ( .I1(n13770), .I2(img[1386]), .O(n25603) );
  ND3S U27272 ( .I1(n26010), .I2(n25604), .I3(n25603), .O(n25605) );
  MUX2 U27273 ( .A(img[1362]), .B(n25605), .S(n29051), .O(n12166) );
  AOI22S U27274 ( .A1(n24415), .A2(img[978]), .B1(n25859), .B2(n30603), .O(
        n25606) );
  ND2S U27275 ( .I1(n26010), .I2(n25606), .O(n25607) );
  AOI22S U27276 ( .A1(n28382), .A2(img[938]), .B1(n13781), .B2(n30604), .O(
        n25608) );
  ND2S U27277 ( .I1(n26010), .I2(n25608), .O(n25609) );
  MUX2 U27278 ( .A(img[978]), .B(n25609), .S(n29145), .O(n12554) );
  AOI22S U27279 ( .A1(n26855), .A2(img[210]), .B1(n28938), .B2(n30605), .O(
        n25610) );
  ND2S U27280 ( .I1(n26010), .I2(n25610), .O(n25611) );
  MUX2 U27281 ( .A(img[170]), .B(n25611), .S(n29148), .O(n13358) );
  AOI22S U27282 ( .A1(n26970), .A2(img[170]), .B1(n25859), .B2(n30606), .O(
        n25612) );
  ND2S U27283 ( .I1(n26010), .I2(n25612), .O(n25613) );
  MUX2 U27284 ( .A(img[210]), .B(n25613), .S(n29151), .O(n13322) );
  AOI22S U27285 ( .A1(n27065), .A2(img[338]), .B1(n13781), .B2(n30607), .O(
        n25614) );
  ND2S U27286 ( .I1(n26010), .I2(n25614), .O(n25615) );
  AOI22S U27287 ( .A1(n27990), .A2(img[298]), .B1(n28343), .B2(n30608), .O(
        n25616) );
  ND2S U27288 ( .I1(n26010), .I2(n25616), .O(n25617) );
  MUX2 U27289 ( .A(img[338]), .B(n25617), .S(n29157), .O(n13190) );
  AOI22S U27290 ( .A1(n26855), .A2(img[466]), .B1(n13781), .B2(n30609), .O(
        n25618) );
  ND2S U27291 ( .I1(n26010), .I2(n25618), .O(n25619) );
  MUX2 U27292 ( .A(img[426]), .B(n25619), .S(n29160), .O(n13102) );
  AOI22S U27293 ( .A1(n25595), .A2(img[426]), .B1(n13781), .B2(n30610), .O(
        n25620) );
  ND2S U27294 ( .I1(n26010), .I2(n25620), .O(n25621) );
  MUX2 U27295 ( .A(img[466]), .B(n25621), .S(n29163), .O(n13066) );
  AOI22S U27296 ( .A1(n27990), .A2(img[1514]), .B1(n29242), .B2(n30611), .O(
        n25622) );
  ND2S U27297 ( .I1(n26010), .I2(n25622), .O(n25623) );
  AOI22S U27298 ( .A1(n25468), .A2(n30612), .B1(n25444), .B2(img[1426]), .O(
        n25625) );
  ND3S U27299 ( .I1(n26010), .I2(n25625), .I3(n25624), .O(n25626) );
  MUX2 U27300 ( .A(img[1514]), .B(n25626), .S(n29099), .O(n12014) );
  AOI22S U27301 ( .A1(n13776), .A2(img[1490]), .B1(n23941), .B2(n30613), .O(
        n25627) );
  ND2S U27302 ( .I1(n26010), .I2(n25627), .O(n25628) );
  AOI22S U27303 ( .A1(n13781), .A2(n30614), .B1(n24946), .B2(img[1450]), .O(
        n25630) );
  ND2S U27304 ( .I1(n13902), .I2(img[1514]), .O(n25629) );
  ND3S U27305 ( .I1(n26010), .I2(n25630), .I3(n25629), .O(n25631) );
  MUX2 U27306 ( .A(n25631), .B(img[1490]), .S(n29091), .O(n12042) );
  AOI22S U27307 ( .A1(n13772), .A2(img[850]), .B1(n25859), .B2(n30615), .O(
        n25632) );
  ND2S U27308 ( .I1(n26010), .I2(n25632), .O(n25633) );
  MUX2 U27309 ( .A(n25633), .B(img[810]), .S(n29166), .O(n12722) );
  INV1S U27310 ( .I(img[850]), .O(n25634) );
  AOI22S U27311 ( .A1(n29435), .A2(img[810]), .B1(n25377), .B2(n25634), .O(
        n25635) );
  ND2S U27312 ( .I1(n13769), .I2(n25635), .O(n25636) );
  AOI22S U27313 ( .A1(n29435), .A2(img[722]), .B1(n25591), .B2(n30616), .O(
        n25637) );
  ND2S U27314 ( .I1(n13769), .I2(n25637), .O(n25638) );
  AOI22S U27315 ( .A1(n13772), .A2(img[682]), .B1(n28695), .B2(n30617), .O(
        n25639) );
  ND2S U27316 ( .I1(n13769), .I2(n25639), .O(n25640) );
  AOI22S U27317 ( .A1(n27685), .A2(img[1130]), .B1(n27511), .B2(n30618), .O(
        n25641) );
  ND2S U27318 ( .I1(n13769), .I2(n25641), .O(n25642) );
  MUX2 U27319 ( .A(n25642), .B(img[1042]), .S(n29122), .O(n12485) );
  AOI22S U27320 ( .A1(n28135), .A2(n30619), .B1(n27919), .B2(img[1042]), .O(
        n25644) );
  ND3S U27321 ( .I1(n26010), .I2(n25644), .I3(n25643), .O(n25645) );
  MUX2 U27322 ( .A(img[1130]), .B(n25645), .S(n29127), .O(n12402) );
  AOI22S U27323 ( .A1(n27065), .A2(img[1106]), .B1(n27511), .B2(n30620), .O(
        n25646) );
  ND2S U27324 ( .I1(n13769), .I2(n25646), .O(n25647) );
  MUX2 U27325 ( .A(n25647), .B(img[1066]), .S(n29115), .O(n12466) );
  AOI22S U27326 ( .A1(n28135), .A2(n30621), .B1(n24313), .B2(img[1066]), .O(
        n25649) );
  ND2S U27327 ( .I1(n13819), .I2(img[1130]), .O(n25648) );
  ND3S U27328 ( .I1(n26010), .I2(n25649), .I3(n25648), .O(n25650) );
  MUX2 U27329 ( .A(img[1106]), .B(n25650), .S(n29119), .O(n12422) );
  AOI22S U27330 ( .A1(n28347), .A2(img[658]), .B1(n28862), .B2(n30622), .O(
        n25651) );
  ND2S U27331 ( .I1(n13769), .I2(n25651), .O(n25652) );
  AOI22S U27332 ( .A1(n13778), .A2(img[746]), .B1(n28162), .B2(n30623), .O(
        n25653) );
  ND2S U27333 ( .I1(n13769), .I2(n25653), .O(n25654) );
  AOI22S U27334 ( .A1(n27110), .A2(img[274]), .B1(n13781), .B2(n30624), .O(
        n25655) );
  ND2S U27335 ( .I1(n13769), .I2(n25655), .O(n25656) );
  MUX2 U27336 ( .A(img[362]), .B(n25656), .S(n29078), .O(n13170) );
  AOI22S U27337 ( .A1(n28347), .A2(img[362]), .B1(n13781), .B2(n30625), .O(
        n25657) );
  ND2S U27338 ( .I1(n13769), .I2(n25657), .O(n25658) );
  AOI22S U27339 ( .A1(n26822), .A2(img[530]), .B1(n13775), .B2(n30626), .O(
        n25659) );
  ND2S U27340 ( .I1(n13769), .I2(n25659), .O(n25660) );
  MUX2 U27341 ( .A(n25660), .B(img[618]), .S(n29024), .O(n12914) );
  AOI22S U27342 ( .A1(n27065), .A2(img[618]), .B1(n29457), .B2(n30627), .O(
        n25661) );
  ND2S U27343 ( .I1(n13769), .I2(n25661), .O(n25662) );
  AOI22S U27344 ( .A1(n29072), .A2(img[18]), .B1(n29457), .B2(n30628), .O(
        n25663) );
  ND2S U27345 ( .I1(n13769), .I2(n25663), .O(n25664) );
  AOI22S U27346 ( .A1(n13777), .A2(img[106]), .B1(n28162), .B2(n30629), .O(
        n25665) );
  ND2S U27347 ( .I1(n13769), .I2(n25665), .O(n25666) );
  MUX2 U27348 ( .A(img[18]), .B(n25666), .S(n29027), .O(n13510) );
  AOI22S U27349 ( .A1(n24415), .A2(img[914]), .B1(n13781), .B2(n30630), .O(
        n25667) );
  ND2S U27350 ( .I1(n13769), .I2(n25667), .O(n25668) );
  AOI22S U27351 ( .A1(n27065), .A2(img[1002]), .B1(n29457), .B2(n30631), .O(
        n25669) );
  ND2S U27352 ( .I1(n13769), .I2(n25669), .O(n25670) );
  MUX2 U27353 ( .A(img[914]), .B(n25670), .S(n29061), .O(n12618) );
  AOI22S U27354 ( .A1(n28347), .A2(img[146]), .B1(n24755), .B2(n30632), .O(
        n25671) );
  ND2S U27355 ( .I1(n13769), .I2(n25671), .O(n25672) );
  MUX2 U27356 ( .A(img[234]), .B(n25672), .S(n29070), .O(n13294) );
  AOI22S U27357 ( .A1(n26101), .A2(img[234]), .B1(n29530), .B2(n30633), .O(
        n25673) );
  ND2S U27358 ( .I1(n13769), .I2(n25673), .O(n25674) );
  MUX2 U27359 ( .A(img[146]), .B(n25674), .S(n29067), .O(n13386) );
  AOI22S U27360 ( .A1(n28382), .A2(img[402]), .B1(n25859), .B2(n30634), .O(
        n25675) );
  ND2S U27361 ( .I1(n13769), .I2(n25675), .O(n25676) );
  MUX2 U27362 ( .A(img[490]), .B(n25676), .S(n29084), .O(n13038) );
  AOI22S U27363 ( .A1(n28347), .A2(img[490]), .B1(n28913), .B2(n30635), .O(
        n25677) );
  ND2S U27364 ( .I1(n13769), .I2(n25677), .O(n25678) );
  INV1S U27365 ( .I(img[874]), .O(n25679) );
  AOI22S U27366 ( .A1(n26970), .A2(img[786]), .B1(n28162), .B2(n25679), .O(
        n25680) );
  ND2S U27367 ( .I1(n13769), .I2(n25680), .O(n25681) );
  AOI22S U27368 ( .A1(n28106), .A2(img[874]), .B1(n25591), .B2(n30636), .O(
        n25682) );
  ND2S U27369 ( .I1(n13769), .I2(n25682), .O(n25683) );
  MUX2 U27370 ( .A(img[786]), .B(n25683), .S(n29102), .O(n12742) );
  AOI22S U27371 ( .A1(n13780), .A2(img[1218]), .B1(n25591), .B2(n30637), .O(
        n25684) );
  ND2S U27372 ( .I1(n13769), .I2(n25684), .O(n25685) );
  MUX2 U27373 ( .A(img[1210]), .B(n25685), .S(n28821), .O(n12318) );
  AOI22S U27374 ( .A1(n28862), .A2(n30638), .B1(n28254), .B2(img[1210]), .O(
        n25687) );
  ND2S U27375 ( .I1(n29124), .I2(img[1274]), .O(n25686) );
  ND3S U27376 ( .I1(n26010), .I2(n25687), .I3(n25686), .O(n25688) );
  MUX2 U27377 ( .A(img[1218]), .B(n25688), .S(n28818), .O(n12314) );
  AOI22S U27378 ( .A1(n13780), .A2(img[1274]), .B1(n28862), .B2(n30639), .O(
        n25689) );
  ND2S U27379 ( .I1(n13769), .I2(n25689), .O(n25690) );
  AOI22S U27380 ( .A1(n29242), .A2(n30640), .B1(n24313), .B2(img[1154]), .O(
        n25692) );
  ND2S U27381 ( .I1(n13820), .I2(img[1218]), .O(n25691) );
  ND3S U27382 ( .I1(n26010), .I2(n25692), .I3(n25691), .O(n25693) );
  MUX2 U27383 ( .A(img[1274]), .B(n25693), .S(n28814), .O(n12254) );
  AOI22S U27384 ( .A1(n13780), .A2(img[2010]), .B1(n28862), .B2(n30641), .O(
        n25694) );
  ND2S U27385 ( .I1(n13769), .I2(n25694), .O(n25695) );
  MUX2 U27386 ( .A(n25695), .B(img[1954]), .S(n28993), .O(n11578) );
  AOI22S U27387 ( .A1(n28037), .A2(n30642), .B1(n24313), .B2(img[1954]), .O(
        n25697) );
  ND2S U27388 ( .I1(n13820), .I2(img[2018]), .O(n25696) );
  ND3S U27389 ( .I1(n26010), .I2(n25697), .I3(n25696), .O(n25698) );
  AOI22S U27390 ( .A1(n13780), .A2(img[2018]), .B1(n29530), .B2(n30643), .O(
        n25699) );
  ND2S U27391 ( .I1(n13769), .I2(n25699), .O(n25700) );
  MUX2 U27392 ( .A(img[1946]), .B(n25700), .S(n29000), .O(n11582) );
  AOI22S U27393 ( .A1(n28037), .A2(n30644), .B1(n25444), .B2(img[1946]), .O(
        n25702) );
  AOI22S U27394 ( .A1(n13899), .A2(img[2010]), .B1(img[2042]), .B2(n13782), 
        .O(n25701) );
  ND3S U27395 ( .I1(n26010), .I2(n25702), .I3(n25701), .O(n25703) );
  MUX2 U27396 ( .A(img[2018]), .B(n25703), .S(n29004), .O(n11514) );
  AOI22S U27397 ( .A1(n28083), .A2(img[1986]), .B1(n13781), .B2(n30645), .O(
        n25704) );
  ND2S U27398 ( .I1(n13769), .I2(n25704), .O(n25705) );
  MUX2 U27399 ( .A(img[1978]), .B(n25705), .S(n29018), .O(n11550) );
  AOI22S U27400 ( .A1(n28037), .A2(n30646), .B1(n24313), .B2(img[1978]), .O(
        n25707) );
  ND3S U27401 ( .I1(n26010), .I2(n25707), .I3(n25706), .O(n25708) );
  MUX2 U27402 ( .A(img[1986]), .B(n25708), .S(n29015), .O(n11546) );
  AOI22S U27403 ( .A1(n28442), .A2(img[2042]), .B1(n29397), .B2(n30647), .O(
        n25709) );
  ND2S U27404 ( .I1(n13769), .I2(n25709), .O(n25710) );
  AOI22S U27405 ( .A1(n28037), .A2(n30648), .B1(n28069), .B2(img[1922]), .O(
        n25712) );
  AOI22S U27406 ( .A1(n13905), .A2(img[1986]), .B1(img[2018]), .B2(n13782), 
        .O(n25711) );
  ND3S U27407 ( .I1(n26010), .I2(n25712), .I3(n25711), .O(n25713) );
  MUX2 U27408 ( .A(img[2042]), .B(n25713), .S(n29011), .O(n11490) );
  AOI22S U27409 ( .A1(n24415), .A2(img[634]), .B1(n28614), .B2(n30649), .O(
        n25714) );
  ND2S U27410 ( .I1(n13769), .I2(n25714), .O(n25715) );
  AOI22S U27411 ( .A1(n28106), .A2(img[514]), .B1(n25591), .B2(n30650), .O(
        n25716) );
  ND2S U27412 ( .I1(n13769), .I2(n25716), .O(n25717) );
  MUX2 U27413 ( .A(n25717), .B(img[634]), .S(n29386), .O(n12898) );
  AOI22S U27414 ( .A1(n27746), .A2(img[1346]), .B1(n25377), .B2(n30651), .O(
        n25718) );
  ND2S U27415 ( .I1(n13769), .I2(n25718), .O(n25719) );
  AOI22S U27416 ( .A1(n28075), .A2(n30652), .B1(n28069), .B2(img[1338]), .O(
        n25721) );
  ND2S U27417 ( .I1(n13905), .I2(img[1402]), .O(n25720) );
  ND3S U27418 ( .I1(n26010), .I2(n25721), .I3(n25720), .O(n25722) );
  MUX2 U27419 ( .A(img[1346]), .B(n25722), .S(n28832), .O(n12182) );
  AOI22S U27420 ( .A1(n29072), .A2(img[1402]), .B1(n28862), .B2(n30653), .O(
        n25723) );
  ND2S U27421 ( .I1(n13769), .I2(n25723), .O(n25724) );
  MUX2 U27422 ( .A(img[1282]), .B(n25724), .S(n28824), .O(n12246) );
  AOI22S U27423 ( .A1(n25062), .A2(n30654), .B1(n28254), .B2(img[1282]), .O(
        n25726) );
  ND3S U27424 ( .I1(n26010), .I2(n25726), .I3(n25725), .O(n25727) );
  MUX2 U27425 ( .A(img[1402]), .B(n25727), .S(n28828), .O(n12130) );
  AOI22S U27426 ( .A1(n29435), .A2(img[250]), .B1(n25859), .B2(n30655), .O(
        n25728) );
  ND2S U27427 ( .I1(n13769), .I2(n25728), .O(n25729) );
  MUX2 U27428 ( .A(n25729), .B(img[130]), .S(n29402), .O(n13402) );
  AOI22S U27429 ( .A1(n25810), .A2(img[130]), .B1(n24374), .B2(n30656), .O(
        n25730) );
  ND2S U27430 ( .I1(n13769), .I2(n25730), .O(n25731) );
  MUX2 U27431 ( .A(img[250]), .B(n25731), .S(n29405), .O(n13277) );
  AOI22S U27432 ( .A1(n25810), .A2(img[378]), .B1(n13775), .B2(n30657), .O(
        n25732) );
  ND2S U27433 ( .I1(n13769), .I2(n25732), .O(n25733) );
  AOI22S U27434 ( .A1(n25810), .A2(img[258]), .B1(n29530), .B2(n30658), .O(
        n25734) );
  ND2S U27435 ( .I1(n13769), .I2(n25734), .O(n25735) );
  MUX2 U27436 ( .A(img[378]), .B(n25735), .S(n29412), .O(n13154) );
  AOI22S U27437 ( .A1(n25810), .A2(img[506]), .B1(n29457), .B2(n30659), .O(
        n25736) );
  ND2S U27438 ( .I1(n13769), .I2(n25736), .O(n25737) );
  MUX2 U27439 ( .A(n25737), .B(img[386]), .S(n29416), .O(n13146) );
  INV1S U27440 ( .I(img[506]), .O(n25738) );
  AOI22S U27441 ( .A1(n13780), .A2(img[386]), .B1(n28862), .B2(n25738), .O(
        n25739) );
  ND2S U27442 ( .I1(n13769), .I2(n25739), .O(n25740) );
  AOI22S U27443 ( .A1(n13780), .A2(img[1474]), .B1(n23941), .B2(n30660), .O(
        n25741) );
  ND2S U27444 ( .I1(n13769), .I2(n25741), .O(n25742) );
  AOI22S U27445 ( .A1(n28075), .A2(n30661), .B1(n28069), .B2(img[1466]), .O(
        n25744) );
  ND2S U27446 ( .I1(n13819), .I2(img[1530]), .O(n25743) );
  ND3S U27447 ( .I1(n26010), .I2(n25744), .I3(n25743), .O(n25745) );
  MUX2 U27448 ( .A(img[1474]), .B(n25745), .S(n28872), .O(n12058) );
  AOI22S U27449 ( .A1(n13780), .A2(img[1530]), .B1(n25591), .B2(n30662), .O(
        n25746) );
  ND2S U27450 ( .I1(n13769), .I2(n25746), .O(n25747) );
  MUX2 U27451 ( .A(img[1410]), .B(n25747), .S(n28864), .O(n12122) );
  AOI22S U27452 ( .A1(n28614), .A2(n30663), .B1(n28254), .B2(img[1410]), .O(
        n25749) );
  ND3S U27453 ( .I1(n26010), .I2(n25749), .I3(n25748), .O(n25750) );
  AOI22S U27454 ( .A1(n13780), .A2(img[890]), .B1(n25591), .B2(n30664), .O(
        n25751) );
  ND2S U27455 ( .I1(n13769), .I2(n25751), .O(n25752) );
  MUX2 U27456 ( .A(img[770]), .B(n25752), .S(n29423), .O(n12758) );
  INV1S U27457 ( .I(img[890]), .O(n25753) );
  AOI22S U27458 ( .A1(n13780), .A2(img[770]), .B1(n29397), .B2(n25753), .O(
        n25754) );
  ND2S U27459 ( .I1(n13769), .I2(n25754), .O(n25755) );
  AOI22S U27460 ( .A1(n13780), .A2(img[762]), .B1(n28913), .B2(n30665), .O(
        n25756) );
  ND2S U27461 ( .I1(n13769), .I2(n25756), .O(n25757) );
  AOI22S U27462 ( .A1(n13780), .A2(img[642]), .B1(n29457), .B2(n30666), .O(
        n25758) );
  ND2S U27463 ( .I1(n13769), .I2(n25758), .O(n25759) );
  AOI22S U27464 ( .A1(n28347), .A2(img[1882]), .B1(n25591), .B2(n30667), .O(
        n25760) );
  ND2S U27465 ( .I1(n13769), .I2(n25760), .O(n25761) );
  AOI22S U27466 ( .A1(n28862), .A2(n30668), .B1(n28069), .B2(img[1826]), .O(
        n25763) );
  ND3S U27467 ( .I1(n26010), .I2(n25763), .I3(n25762), .O(n25764) );
  MUX2 U27468 ( .A(img[1882]), .B(n25764), .S(n28896), .O(n11650) );
  AOI22S U27469 ( .A1(n29072), .A2(img[1890]), .B1(n27049), .B2(n30669), .O(
        n25765) );
  ND2S U27470 ( .I1(n13769), .I2(n25765), .O(n25766) );
  AOI22S U27471 ( .A1(n28862), .A2(n30670), .B1(n28254), .B2(img[1818]), .O(
        n25768) );
  AOI22S U27472 ( .A1(n13905), .A2(img[1882]), .B1(img[1914]), .B2(n13782), 
        .O(n25767) );
  ND3S U27473 ( .I1(n26010), .I2(n25768), .I3(n25767), .O(n25769) );
  MUX2 U27474 ( .A(img[1890]), .B(n25769), .S(n28903), .O(n11638) );
  AOI22S U27475 ( .A1(n26822), .A2(img[1858]), .B1(n27049), .B2(n30671), .O(
        n25770) );
  ND2S U27476 ( .I1(n13769), .I2(n25770), .O(n25771) );
  MUX2 U27477 ( .A(img[1850]), .B(n25771), .S(n28919), .O(n11682) );
  AOI22S U27478 ( .A1(n28343), .A2(n30672), .B1(n28254), .B2(img[1850]), .O(
        n25773) );
  ND3S U27479 ( .I1(n26010), .I2(n25773), .I3(n25772), .O(n25774) );
  MUX2 U27480 ( .A(img[1858]), .B(n25774), .S(n28916), .O(n11670) );
  AOI22S U27481 ( .A1(n29435), .A2(img[1914]), .B1(n27049), .B2(n30673), .O(
        n25775) );
  ND2S U27482 ( .I1(n13769), .I2(n25775), .O(n25776) );
  AOI22S U27483 ( .A1(n28592), .A2(n30674), .B1(n28254), .B2(img[1794]), .O(
        n257780) );
  AOI22S U27484 ( .A1(n13905), .A2(img[1858]), .B1(img[1890]), .B2(n13782), 
        .O(n257770) );
  ND3S U27485 ( .I1(n26010), .I2(n257780), .I3(n257770), .O(n25779) );
  MUX2 U27486 ( .A(img[1914]), .B(n25779), .S(n28911), .O(n11618) );
  AOI22S U27487 ( .A1(n25810), .A2(img[1754]), .B1(n27049), .B2(n30675), .O(
        n25780) );
  ND2S U27488 ( .I1(n26010), .I2(n25780), .O(n25781) );
  AOI22S U27489 ( .A1(n28862), .A2(n30676), .B1(n28069), .B2(img[1698]), .O(
        n25783) );
  ND2S U27490 ( .I1(n13820), .I2(img[1762]), .O(n25782) );
  ND3S U27491 ( .I1(n26010), .I2(n25783), .I3(n25782), .O(n25784) );
  MUX2 U27492 ( .A(img[1754]), .B(n25784), .S(n28926), .O(n11774) );
  AOI22S U27493 ( .A1(n25810), .A2(img[1762]), .B1(n27049), .B2(n30677), .O(
        n25785) );
  ND2S U27494 ( .I1(n26010), .I2(n25785), .O(n25786) );
  AOI22S U27495 ( .A1(n25591), .A2(n30678), .B1(n28069), .B2(img[1690]), .O(
        n25788) );
  AOI22S U27496 ( .A1(n13905), .A2(img[1754]), .B1(img[1786]), .B2(n13782), 
        .O(n25787) );
  ND3S U27497 ( .I1(n26010), .I2(n25788), .I3(n25787), .O(n25789) );
  MUX2 U27498 ( .A(img[1762]), .B(n25789), .S(n28933), .O(n11770) );
  AOI22S U27499 ( .A1(n25810), .A2(img[1730]), .B1(n29397), .B2(n30679), .O(
        n25790) );
  ND2S U27500 ( .I1(n26010), .I2(n25790), .O(n25791) );
  AOI22S U27501 ( .A1(n29096), .A2(n30680), .B1(n28069), .B2(img[1722]), .O(
        n25793) );
  ND3S U27502 ( .I1(n26010), .I2(n25793), .I3(n25792), .O(n25794) );
  MUX2 U27503 ( .A(img[1730]), .B(n25794), .S(n28945), .O(n11802) );
  AOI22S U27504 ( .A1(n25810), .A2(img[1786]), .B1(n27049), .B2(n30681), .O(
        n25795) );
  ND2S U27505 ( .I1(n26010), .I2(n25795), .O(n25796) );
  AOI22S U27506 ( .A1(n28938), .A2(n30682), .B1(n28069), .B2(img[1666]), .O(
        n25798) );
  AOI22S U27507 ( .A1(n13905), .A2(img[1730]), .B1(img[1762]), .B2(n13782), 
        .O(n25797) );
  ND3S U27508 ( .I1(n26010), .I2(n25798), .I3(n25797), .O(n25799) );
  MUX2 U27509 ( .A(img[1786]), .B(n25799), .S(n28941), .O(n11742) );
  AOI22S U27510 ( .A1(n25810), .A2(img[1626]), .B1(n27049), .B2(n30683), .O(
        n25800) );
  ND2S U27511 ( .I1(n26010), .I2(n25800), .O(n25801) );
  AOI22S U27512 ( .A1(n13781), .A2(n30684), .B1(n24946), .B2(img[1570]), .O(
        n25803) );
  ND3S U27513 ( .I1(n26010), .I2(n25803), .I3(n25802), .O(n25804) );
  MUX2 U27514 ( .A(img[1626]), .B(n25804), .S(n28955), .O(n11906) );
  AOI22S U27515 ( .A1(n25810), .A2(img[1634]), .B1(n27049), .B2(n30685), .O(
        n25805) );
  ND2S U27516 ( .I1(n26010), .I2(n25805), .O(n25806) );
  AOI22S U27517 ( .A1(n28037), .A2(n30686), .B1(n28069), .B2(img[1562]), .O(
        n25808) );
  AOI22S U27518 ( .A1(n13903), .A2(img[1626]), .B1(img[1658]), .B2(n13782), 
        .O(n25807) );
  ND3S U27519 ( .I1(n26010), .I2(n25808), .I3(n25807), .O(n25809) );
  MUX2 U27520 ( .A(img[1634]), .B(n25809), .S(n28962), .O(n11893) );
  AOI22S U27521 ( .A1(n25810), .A2(img[1602]), .B1(n27049), .B2(n30687), .O(
        n25811) );
  ND2S U27522 ( .I1(n26010), .I2(n25811), .O(n25812) );
  AOI22S U27523 ( .A1(n25468), .A2(n30688), .B1(n28069), .B2(img[1594]), .O(
        n25814) );
  ND2S U27524 ( .I1(n13770), .I2(img[1658]), .O(n25813) );
  ND3S U27525 ( .I1(n26010), .I2(n25814), .I3(n25813), .O(n25815) );
  MUX2 U27526 ( .A(img[1602]), .B(n25815), .S(n28973), .O(n11926) );
  AOI22S U27527 ( .A1(n29072), .A2(img[1658]), .B1(n24374), .B2(n30689), .O(
        n25816) );
  ND2S U27528 ( .I1(n26010), .I2(n25816), .O(n25817) );
  AOI22S U27529 ( .A1(n28162), .A2(n30690), .B1(n24313), .B2(img[1538]), .O(
        n25819) );
  AOI22S U27530 ( .A1(n13899), .A2(img[1602]), .B1(img[1634]), .B2(n13782), 
        .O(n25818) );
  ND3S U27531 ( .I1(n26010), .I2(n25819), .I3(n25818), .O(n25820) );
  MUX2 U27532 ( .A(img[1658]), .B(n25820), .S(n28969), .O(n11874) );
  AOI22S U27533 ( .A1(n25810), .A2(img[1090]), .B1(n23941), .B2(n30691), .O(
        n25821) );
  ND2S U27534 ( .I1(n26010), .I2(n25821), .O(n25822) );
  AOI22S U27535 ( .A1(n28614), .A2(n30692), .B1(n24313), .B2(img[1082]), .O(
        n25824) );
  ND3S U27536 ( .I1(n26010), .I2(n25824), .I3(n25823), .O(n25825) );
  MUX2 U27537 ( .A(img[1090]), .B(n25825), .S(n28987), .O(n12442) );
  AOI22S U27538 ( .A1(n28347), .A2(img[1146]), .B1(n28913), .B2(n30693), .O(
        n25826) );
  ND2S U27539 ( .I1(n26010), .I2(n25826), .O(n25827) );
  AOI22S U27540 ( .A1(n25591), .A2(n30694), .B1(n24313), .B2(img[1026]), .O(
        n25829) );
  ND2S U27541 ( .I1(n13905), .I2(img[1090]), .O(n25828) );
  ND3S U27542 ( .I1(n26010), .I2(n25829), .I3(n25828), .O(n25830) );
  MUX2 U27543 ( .A(img[1146]), .B(n25830), .S(n28983), .O(n12386) );
  AOI22S U27544 ( .A1(n27746), .A2(img[122]), .B1(n13775), .B2(n30695), .O(
        n25831) );
  ND2S U27545 ( .I1(n26010), .I2(n25831), .O(n25832) );
  AOI22S U27546 ( .A1(n13776), .A2(img[2]), .B1(n23941), .B2(n30696), .O(
        n25833) );
  ND2S U27547 ( .I1(n26010), .I2(n25833), .O(n25834) );
  MUX2 U27548 ( .A(img[122]), .B(n25834), .S(n29392), .O(n13410) );
  AOI22S U27549 ( .A1(n28347), .A2(img[1018]), .B1(n28862), .B2(n30697), .O(
        n25835) );
  ND2S U27550 ( .I1(n26010), .I2(n25835), .O(n25836) );
  AOI22S U27551 ( .A1(n28106), .A2(img[898]), .B1(n29397), .B2(n30698), .O(
        n25837) );
  ND2S U27552 ( .I1(n26010), .I2(n25837), .O(n25838) );
  MUX2 U27553 ( .A(img[1018]), .B(n25838), .S(n29399), .O(n12510) );
  AOI22S U27554 ( .A1(n27065), .A2(img[586]), .B1(n13775), .B2(n30699), .O(
        n25839) );
  ND2S U27555 ( .I1(n26010), .I2(n25839), .O(n25840) );
  MUX2 U27556 ( .A(n25840), .B(img[562]), .S(n28578), .O(n12966) );
  AOI22S U27557 ( .A1(n28347), .A2(img[562]), .B1(n13775), .B2(n30700), .O(
        n25841) );
  ND2S U27558 ( .I1(n26010), .I2(n25841), .O(n25842) );
  MUX2 U27559 ( .A(n25842), .B(img[586]), .S(n28581), .O(n12946) );
  AOI22S U27560 ( .A1(n28347), .A2(img[74]), .B1(n25859), .B2(n30701), .O(
        n25843) );
  ND2S U27561 ( .I1(n26010), .I2(n25843), .O(n25844) );
  MUX2 U27562 ( .A(img[50]), .B(n25844), .S(n28584), .O(n13483) );
  AOI22S U27563 ( .A1(n28442), .A2(img[50]), .B1(n25859), .B2(n30702), .O(
        n25845) );
  ND2S U27564 ( .I1(n26010), .I2(n25845), .O(n25846) );
  AOI22S U27565 ( .A1(n28840), .A2(img[970]), .B1(n25859), .B2(n30703), .O(
        n25847) );
  ND2S U27566 ( .I1(n26010), .I2(n25847), .O(n25848) );
  AOI22S U27567 ( .A1(n27065), .A2(img[946]), .B1(n25859), .B2(n30704), .O(
        n25849) );
  ND2S U27568 ( .I1(n26010), .I2(n25849), .O(n25850) );
  MUX2 U27569 ( .A(img[970]), .B(n25850), .S(n28623), .O(n12558) );
  AOI22S U27570 ( .A1(n26101), .A2(img[202]), .B1(n25859), .B2(n30705), .O(
        n25851) );
  ND2S U27571 ( .I1(n26010), .I2(n25851), .O(n25852) );
  MUX2 U27572 ( .A(img[178]), .B(n25852), .S(n28626), .O(n13354) );
  AOI22S U27573 ( .A1(n26855), .A2(img[178]), .B1(n25859), .B2(n30706), .O(
        n25853) );
  ND2S U27574 ( .I1(n26010), .I2(n25853), .O(n25854) );
  MUX2 U27575 ( .A(img[202]), .B(n25854), .S(n28629), .O(n13326) );
  AOI22S U27576 ( .A1(n25595), .A2(img[458]), .B1(n25859), .B2(n30707), .O(
        n25855) );
  ND2S U27577 ( .I1(n26010), .I2(n25855), .O(n25856) );
  AOI22S U27578 ( .A1(n26101), .A2(img[434]), .B1(n25859), .B2(n30708), .O(
        n25857) );
  ND2S U27579 ( .I1(n26010), .I2(n25857), .O(n25858) );
  MUX2 U27580 ( .A(n25858), .B(img[458]), .S(n28641), .O(n13070) );
  AOI22S U27581 ( .A1(n13780), .A2(img[842]), .B1(n25859), .B2(n30709), .O(
        n25860) );
  ND2S U27582 ( .I1(n26010), .I2(n25860), .O(n25861) );
  INV1S U27583 ( .I(img[842]), .O(n25862) );
  AOI22S U27584 ( .A1(n25595), .A2(img[818]), .B1(n27049), .B2(n25862), .O(
        n25863) );
  ND2S U27585 ( .I1(n26010), .I2(n25863), .O(n25864) );
  AOI22S U27586 ( .A1(n28347), .A2(img[330]), .B1(n24755), .B2(n30710), .O(
        n25865) );
  ND2S U27587 ( .I1(n26010), .I2(n25865), .O(n25866) );
  MUX2 U27588 ( .A(img[306]), .B(n25866), .S(n28632), .O(n13222) );
  AOI22S U27589 ( .A1(n28106), .A2(img[306]), .B1(n29530), .B2(n30711), .O(
        n25867) );
  ND2S U27590 ( .I1(n26010), .I2(n25867), .O(n25868) );
  AOI22S U27591 ( .A1(n28083), .A2(img[714]), .B1(n24193), .B2(n30712), .O(
        n25869) );
  ND2S U27592 ( .I1(n26010), .I2(n25869), .O(n25870) );
  AOI22S U27593 ( .A1(n25595), .A2(img[690]), .B1(n24374), .B2(n30713), .O(
        n25871) );
  ND2S U27594 ( .I1(n26010), .I2(n25871), .O(n25872) );
  AOI22S U27595 ( .A1(n27065), .A2(img[90]), .B1(n25377), .B2(n30714), .O(
        n25873) );
  ND2S U27596 ( .I1(n26010), .I2(n25873), .O(n25874) );
  AOI22S U27597 ( .A1(n24415), .A2(img[34]), .B1(n29457), .B2(n30715), .O(
        n25875) );
  ND2S U27598 ( .I1(n26010), .I2(n25875), .O(n25876) );
  MUX2 U27599 ( .A(img[90]), .B(n25876), .S(n29339), .O(n13442) );
  AOI22S U27600 ( .A1(n29414), .A2(img[1250]), .B1(n13781), .B2(n30716), .O(
        n25877) );
  ND2S U27601 ( .I1(n26010), .I2(n25877), .O(n25878) );
  AOI22S U27602 ( .A1(n28135), .A2(n30717), .B1(n28069), .B2(img[1178]), .O(
        n25880) );
  ND2S U27603 ( .I1(n13770), .I2(img[1242]), .O(n25879) );
  ND3S U27604 ( .I1(n26010), .I2(n25880), .I3(n25879), .O(n25881) );
  MUX2 U27605 ( .A(img[1250]), .B(n25881), .S(n29218), .O(n12282) );
  AOI22S U27606 ( .A1(n26822), .A2(img[1242]), .B1(n29407), .B2(n30718), .O(
        n25882) );
  ND2S U27607 ( .I1(n26010), .I2(n25882), .O(n25883) );
  MUX2 U27608 ( .A(n25883), .B(img[1186]), .S(n29207), .O(n12346) );
  AOI22S U27609 ( .A1(n27049), .A2(n30719), .B1(n28069), .B2(img[1186]), .O(
        n25885) );
  ND2S U27610 ( .I1(n13770), .I2(img[1250]), .O(n25884) );
  ND3S U27611 ( .I1(n26010), .I2(n25885), .I3(n25884), .O(n25886) );
  MUX2 U27612 ( .A(img[1242]), .B(n25886), .S(n29211), .O(n12286) );
  AOI22S U27613 ( .A1(n27722), .A2(img[1378]), .B1(n29457), .B2(n30720), .O(
        n25887) );
  ND2S U27614 ( .I1(n26010), .I2(n25887), .O(n25888) );
  MUX2 U27615 ( .A(img[1306]), .B(n25888), .S(n29240), .O(n12226) );
  AOI22S U27616 ( .A1(n28182), .A2(n30721), .B1(n28069), .B2(img[1306]), .O(
        n25890) );
  ND3S U27617 ( .I1(n26010), .I2(n25890), .I3(n25889), .O(n25891) );
  MUX2 U27618 ( .A(img[1378]), .B(n25891), .S(n29245), .O(n12150) );
  AOI22S U27619 ( .A1(n13780), .A2(img[1370]), .B1(n24193), .B2(n30722), .O(
        n25892) );
  ND2S U27620 ( .I1(n26010), .I2(n25892), .O(n25893) );
  MUX2 U27621 ( .A(n25893), .B(img[1314]), .S(n29233), .O(n12214) );
  AOI22S U27622 ( .A1(n29194), .A2(n30723), .B1(n26091), .B2(img[1314]), .O(
        n25895) );
  ND2S U27623 ( .I1(n13770), .I2(img[1378]), .O(n258940) );
  ND3S U27624 ( .I1(n26010), .I2(n25895), .I3(n258940), .O(n25896) );
  MUX2 U27625 ( .A(img[1370]), .B(n25896), .S(n29237), .O(n12162) );
  AOI22S U27626 ( .A1(n27957), .A2(img[218]), .B1(n24374), .B2(n30724), .O(
        n25897) );
  ND2S U27627 ( .I1(n26010), .I2(n25897), .O(n25898) );
  MUX2 U27628 ( .A(img[162]), .B(n25898), .S(n29355), .O(n13370) );
  AOI22S U27629 ( .A1(n29435), .A2(img[162]), .B1(n13775), .B2(n30725), .O(
        n25899) );
  ND2S U27630 ( .I1(n26010), .I2(n25899), .O(n25900) );
  MUX2 U27631 ( .A(img[218]), .B(n25900), .S(n29351), .O(n13310) );
  AOI22S U27632 ( .A1(n29072), .A2(img[346]), .B1(n13779), .B2(n30726), .O(
        n25901) );
  ND2S U27633 ( .I1(n26010), .I2(n25901), .O(n25902) );
  AOI22S U27634 ( .A1(n27722), .A2(img[290]), .B1(n13779), .B2(n30727), .O(
        n25904) );
  ND2S U27635 ( .I1(n13769), .I2(n25904), .O(n25905) );
  MUX2 U27636 ( .A(img[346]), .B(n25905), .S(n29358), .O(n13186) );
  AOI22S U27637 ( .A1(n13772), .A2(img[474]), .B1(n13779), .B2(n30728), .O(
        n25906) );
  ND2S U27638 ( .I1(n13769), .I2(n25906), .O(n25907) );
  AOI22S U27639 ( .A1(n13772), .A2(img[418]), .B1(n13779), .B2(n30729), .O(
        n25908) );
  ND2S U27640 ( .I1(n13769), .I2(n25908), .O(n25909) );
  MUX2 U27641 ( .A(img[474]), .B(n25909), .S(n29364), .O(n13054) );
  AOI22S U27642 ( .A1(n13772), .A2(img[1506]), .B1(n13779), .B2(n30730), .O(
        n25910) );
  ND2S U27643 ( .I1(n13769), .I2(n25910), .O(n25911) );
  MUX2 U27644 ( .A(n25911), .B(img[1434]), .S(n29255), .O(n12094) );
  AOI22S U27645 ( .A1(n28075), .A2(n30731), .B1(n26091), .B2(img[1434]), .O(
        n25913) );
  ND3S U27646 ( .I1(n26010), .I2(n25913), .I3(n25912), .O(n25914) );
  MUX2 U27647 ( .A(img[1506]), .B(n25914), .S(n29261), .O(n12026) );
  AOI22S U27648 ( .A1(n13772), .A2(img[1498]), .B1(n28862), .B2(n30732), .O(
        n25915) );
  ND2S U27649 ( .I1(n13769), .I2(n25915), .O(n25916) );
  MUX2 U27650 ( .A(n25916), .B(img[1442]), .S(n29248), .O(n12090) );
  AOI22S U27651 ( .A1(n28037), .A2(n30733), .B1(n26091), .B2(img[1442]), .O(
        n25918) );
  ND3S U27652 ( .I1(n26010), .I2(n25918), .I3(n25917), .O(n25919) );
  AOI22S U27653 ( .A1(n27065), .A2(img[858]), .B1(n13781), .B2(n30734), .O(
        n25920) );
  ND2S U27654 ( .I1(n13769), .I2(n25920), .O(n25921) );
  MUX2 U27655 ( .A(n25921), .B(img[802]), .S(n29374), .O(n12726) );
  INV1S U27656 ( .I(img[858]), .O(n25922) );
  AOI22S U27657 ( .A1(n13777), .A2(img[802]), .B1(n24755), .B2(n25922), .O(
        n25923) );
  ND2S U27658 ( .I1(n13769), .I2(n25923), .O(n25924) );
  AOI22S U27659 ( .A1(n25810), .A2(img[730]), .B1(n28862), .B2(n30735), .O(
        n25925) );
  ND2S U27660 ( .I1(n13769), .I2(n25925), .O(n25926) );
  AOI22S U27661 ( .A1(n28347), .A2(img[674]), .B1(n29530), .B2(n30736), .O(
        n25927) );
  ND2S U27662 ( .I1(n13769), .I2(n25927), .O(n25928) );
  AOI22S U27663 ( .A1(n28347), .A2(img[1122]), .B1(n24755), .B2(n30737), .O(
        n25929) );
  ND2S U27664 ( .I1(n13769), .I2(n25929), .O(n25930) );
  AOI22S U27665 ( .A1(n28037), .A2(n30738), .B1(n26091), .B2(img[1050]), .O(
        n25932) );
  ND3S U27666 ( .I1(n26010), .I2(n25932), .I3(n25931), .O(n25933) );
  MUX2 U27667 ( .A(img[1122]), .B(n25933), .S(n29198), .O(n12406) );
  AOI22S U27668 ( .A1(n25810), .A2(img[1114]), .B1(n28433), .B2(n30739), .O(
        n25934) );
  ND2S U27669 ( .I1(n13769), .I2(n25934), .O(n25935) );
  MUX2 U27670 ( .A(n25935), .B(img[1058]), .S(n29185), .O(n12470) );
  AOI22S U27671 ( .A1(n28075), .A2(n30740), .B1(n26091), .B2(img[1058]), .O(
        n25937) );
  ND3S U27672 ( .I1(n26010), .I2(n25937), .I3(n25936), .O(n25938) );
  MUX2 U27673 ( .A(img[1114]), .B(n25938), .S(n29189), .O(n12418) );
  AOI22S U27674 ( .A1(n28106), .A2(img[602]), .B1(n13781), .B2(n30741), .O(
        n25939) );
  ND2S U27675 ( .I1(n13769), .I2(n25939), .O(n25940) );
  MUX2 U27676 ( .A(n25940), .B(img[546]), .S(n29481), .O(n12986) );
  AOI22S U27677 ( .A1(n27990), .A2(img[546]), .B1(n28343), .B2(n30742), .O(
        n25941) );
  ND2S U27678 ( .I1(n13769), .I2(n25941), .O(n25942) );
  MUX2 U27679 ( .A(n25942), .B(img[602]), .S(n29478), .O(n12930) );
  AOI22S U27680 ( .A1(n27990), .A2(img[986]), .B1(n29530), .B2(n30743), .O(
        n25943) );
  ND2S U27681 ( .I1(n13769), .I2(n25943), .O(n25944) );
  MUX2 U27682 ( .A(n25944), .B(img[930]), .S(n29348), .O(n12602) );
  AOI22S U27683 ( .A1(n27990), .A2(img[930]), .B1(n13781), .B2(n30744), .O(
        n25945) );
  ND2S U27684 ( .I1(n13769), .I2(n25945), .O(n25946) );
  AOI22S U27685 ( .A1(n27990), .A2(img[538]), .B1(n27049), .B2(n30745), .O(
        n25947) );
  ND2S U27686 ( .I1(n13769), .I2(n25947), .O(n25948) );
  MUX2 U27687 ( .A(n25948), .B(img[610]), .S(n29286), .O(n12918) );
  AOI22S U27688 ( .A1(n13772), .A2(img[610]), .B1(n13779), .B2(n30746), .O(
        n25949) );
  ND2S U27689 ( .I1(n13769), .I2(n25949), .O(n25950) );
  AOI22S U27690 ( .A1(n13772), .A2(img[26]), .B1(n13781), .B2(n30747), .O(
        n25951) );
  ND2S U27691 ( .I1(n13769), .I2(n25951), .O(n25952) );
  MUX2 U27692 ( .A(img[98]), .B(n25952), .S(n29280), .O(n13430) );
  AOI22S U27693 ( .A1(n13772), .A2(img[98]), .B1(n29530), .B2(n30748), .O(
        n25953) );
  ND2S U27694 ( .I1(n13769), .I2(n25953), .O(n25954) );
  AOI22S U27695 ( .A1(n13772), .A2(img[922]), .B1(n27049), .B2(n30749), .O(
        n25955) );
  ND2S U27696 ( .I1(n13769), .I2(n25955), .O(n25956) );
  MUX2 U27697 ( .A(img[994]), .B(n25956), .S(n29224), .O(n12538) );
  AOI22S U27698 ( .A1(n13772), .A2(img[994]), .B1(n29530), .B2(n30750), .O(
        n25957) );
  ND2S U27699 ( .I1(n13769), .I2(n25957), .O(n25958) );
  AOI22S U27700 ( .A1(n13772), .A2(img[154]), .B1(n29242), .B2(n30751), .O(
        n25959) );
  ND2S U27701 ( .I1(n13769), .I2(n25959), .O(n25960) );
  MUX2 U27702 ( .A(img[226]), .B(n25960), .S(n29267), .O(n13306) );
  AOI22S U27703 ( .A1(n13772), .A2(img[226]), .B1(n28162), .B2(n30752), .O(
        n25961) );
  ND2S U27704 ( .I1(n13769), .I2(n25961), .O(n25962) );
  MUX2 U27705 ( .A(img[154]), .B(n25962), .S(n29264), .O(n13374) );
  AOI22S U27706 ( .A1(n28347), .A2(img[282]), .B1(n25859), .B2(n30753), .O(
        n25963) );
  ND2S U27707 ( .I1(n13769), .I2(n25963), .O(n25964) );
  MUX2 U27708 ( .A(img[354]), .B(n25964), .S(n29182), .O(n13174) );
  AOI22S U27709 ( .A1(n26101), .A2(img[354]), .B1(n13781), .B2(n30754), .O(
        n25965) );
  ND2S U27710 ( .I1(n13769), .I2(n25965), .O(n25966) );
  AOI22S U27711 ( .A1(n13772), .A2(img[410]), .B1(n13781), .B2(n30755), .O(
        n25967) );
  ND2S U27712 ( .I1(n13769), .I2(n25967), .O(n25968) );
  MUX2 U27713 ( .A(img[482]), .B(n25968), .S(n29273), .O(n13050) );
  AOI22S U27714 ( .A1(n25595), .A2(img[482]), .B1(n13781), .B2(n30756), .O(
        n25969) );
  ND2S U27715 ( .I1(n26010), .I2(n25969), .O(n25970) );
  AOI22S U27716 ( .A1(n27990), .A2(img[794]), .B1(n13781), .B2(n30757), .O(
        n25971) );
  ND2S U27717 ( .I1(n26010), .I2(n25971), .O(n25972) );
  AOI22S U27718 ( .A1(n27990), .A2(img[866]), .B1(n28182), .B2(n30758), .O(
        n25973) );
  ND2S U27719 ( .I1(n26010), .I2(n25973), .O(n25974) );
  MUX2 U27720 ( .A(img[794]), .B(n25974), .S(n29227), .O(n12738) );
  AOI22S U27721 ( .A1(n27990), .A2(img[666]), .B1(n28614), .B2(n30759), .O(
        n25975) );
  ND2S U27722 ( .I1(n26010), .I2(n25975), .O(n25976) );
  AOI22S U27723 ( .A1(n27990), .A2(img[738]), .B1(n28162), .B2(n30760), .O(
        n25977) );
  ND2S U27724 ( .I1(n26010), .I2(n25977), .O(n25978) );
  AOI22S U27725 ( .A1(n27990), .A2(img[570]), .B1(n28862), .B2(n30761), .O(
        n25979) );
  ND2S U27726 ( .I1(n26010), .I2(n25979), .O(n25980) );
  MUX2 U27727 ( .A(n25980), .B(img[578]), .S(n28799), .O(n12950) );
  AOI22S U27728 ( .A1(n27990), .A2(img[66]), .B1(n27511), .B2(n30762), .O(
        n25981) );
  ND2S U27729 ( .I1(n26010), .I2(n25981), .O(n25982) );
  AOI22S U27730 ( .A1(n27990), .A2(img[58]), .B1(n25062), .B2(n30763), .O(
        n25983) );
  ND2S U27731 ( .I1(n26010), .I2(n25983), .O(n25984) );
  MUX2 U27732 ( .A(img[66]), .B(n25984), .S(n28804), .O(n13462) );
  AOI22S U27733 ( .A1(n28382), .A2(img[962]), .B1(n29407), .B2(n30764), .O(
        n25985) );
  ND2S U27734 ( .I1(n26010), .I2(n25985), .O(n25986) );
  MUX2 U27735 ( .A(img[954]), .B(n25986), .S(n28842), .O(n12574) );
  AOI22S U27736 ( .A1(n28382), .A2(img[954]), .B1(n24755), .B2(n30765), .O(
        n25987) );
  ND2S U27737 ( .I1(n26010), .I2(n25987), .O(n25988) );
  AOI22S U27738 ( .A1(n28382), .A2(img[194]), .B1(n23918), .B2(n30766), .O(
        n25989) );
  ND2S U27739 ( .I1(n26010), .I2(n25989), .O(n25990) );
  MUX2 U27740 ( .A(img[186]), .B(n25990), .S(n28848), .O(n13342) );
  AOI22S U27741 ( .A1(n28382), .A2(img[186]), .B1(n25062), .B2(n30767), .O(
        n25991) );
  ND2S U27742 ( .I1(n26010), .I2(n25991), .O(n25992) );
  MUX2 U27743 ( .A(img[194]), .B(n25992), .S(n28845), .O(n13338) );
  AOI22S U27744 ( .A1(n29129), .A2(img[322]), .B1(n27735), .B2(n30768), .O(
        n25993) );
  ND2S U27745 ( .I1(n26010), .I2(n25993), .O(n25994) );
  AOI22S U27746 ( .A1(n26855), .A2(img[314]), .B1(n25062), .B2(n30769), .O(
        n25995) );
  ND2S U27747 ( .I1(n26010), .I2(n25995), .O(n25996) );
  MUX2 U27748 ( .A(img[322]), .B(n25996), .S(n28851), .O(n13206) );
  AOI22S U27749 ( .A1(n24415), .A2(img[450]), .B1(n25591), .B2(n30770), .O(
        n25997) );
  ND2S U27750 ( .I1(n26010), .I2(n25997), .O(n25998) );
  AOI22S U27751 ( .A1(n26101), .A2(img[442]), .B1(n28343), .B2(n30771), .O(
        n25999) );
  ND2S U27752 ( .I1(n26010), .I2(n25999), .O(n26000) );
  INV1S U27753 ( .I(img[826]), .O(n26001) );
  AOI22S U27754 ( .A1(n29129), .A2(img[834]), .B1(n25591), .B2(n26001), .O(
        n26002) );
  ND2S U27755 ( .I1(n26010), .I2(n26002), .O(n26003) );
  INV1S U27756 ( .I(img[834]), .O(n26004) );
  AOI22S U27757 ( .A1(n27990), .A2(img[826]), .B1(n25062), .B2(n26004), .O(
        n26005) );
  ND2S U27758 ( .I1(n26010), .I2(n26005), .O(n26006) );
  MUX2 U27759 ( .A(n26006), .B(img[834]), .S(n28879), .O(n12694) );
  AOI22S U27760 ( .A1(n28643), .A2(img[706]), .B1(n29194), .B2(n30772), .O(
        n26007) );
  ND2S U27761 ( .I1(n26010), .I2(n26007), .O(n26008) );
  AOI22S U27762 ( .A1(n26101), .A2(img[698]), .B1(n28913), .B2(n30773), .O(
        n26009) );
  ND2S U27763 ( .I1(n26010), .I2(n26009), .O(n26011) );
  OAI22S U27764 ( .A1(n26013), .A2(n28530), .B1(n13897), .B2(n26012), .O(
        n26014) );
  AOI12HS U27765 ( .B1(n28534), .B2(n26015), .A1(n26014), .O(n26016) );
  ND2S U27766 ( .I1(n28550), .I2(A67_shift[77]), .O(n26018) );
  AOI22S U27767 ( .A1(n28554), .A2(A67_shift[109]), .B1(n28551), .B2(
        A67_shift[205]), .O(n26017) );
  NR2 U27768 ( .I1(n26020), .I2(n26019), .O(n26023) );
  AOI22S U27769 ( .A1(n28546), .A2(A67_shift[173]), .B1(n28545), .B2(
        A67_shift[45]), .O(n26021) );
  ND2S U27770 ( .I1(n28550), .I2(A67_shift[93]), .O(n26025) );
  AOI22S U27771 ( .A1(n28554), .A2(A67_shift[125]), .B1(n28551), .B2(
        A67_shift[221]), .O(n26024) );
  NR2 U27772 ( .I1(n26027), .I2(n26026), .O(n26030) );
  AOI22S U27773 ( .A1(n28546), .A2(A67_shift[189]), .B1(n28545), .B2(
        A67_shift[61]), .O(n26028) );
  ND2S U27774 ( .I1(n28564), .I2(gray_avg_out[5]), .O(n26035) );
  ND2S U27775 ( .I1(n28565), .I2(gray_weight_out[5]), .O(n26034) );
  ND2S U27776 ( .I1(n28566), .I2(gray_max_out[5]), .O(n26033) );
  AOI22S U27777 ( .A1(n26101), .A2(img[613]), .B1(n28135), .B2(n30774), .O(
        n26040) );
  ND2S U27778 ( .I1(n26534), .I2(n26040), .O(n26041) );
  MUX2 U27779 ( .A(img[541]), .B(n26041), .S(n29283), .O(n12991) );
  AOI22S U27780 ( .A1(n26101), .A2(img[541]), .B1(n13775), .B2(n30775), .O(
        n26042) );
  ND2S U27781 ( .I1(n26534), .I2(n26042), .O(n26043) );
  MUX2 U27782 ( .A(n26043), .B(img[613]), .S(n29286), .O(n12921) );
  AOI22S U27783 ( .A1(n26101), .A2(img[101]), .B1(n27735), .B2(n30776), .O(
        n26044) );
  ND2S U27784 ( .I1(n26534), .I2(n26044), .O(n26045) );
  MUX2 U27785 ( .A(img[29]), .B(n26045), .S(n29276), .O(n13503) );
  AOI22S U27786 ( .A1(n28382), .A2(img[29]), .B1(n27511), .B2(n30777), .O(
        n26046) );
  ND2S U27787 ( .I1(n26534), .I2(n26046), .O(n26047) );
  MUX2 U27788 ( .A(img[101]), .B(n26047), .S(n29280), .O(n13433) );
  AOI22S U27789 ( .A1(n28382), .A2(img[1245]), .B1(n24193), .B2(n30778), .O(
        n26048) );
  ND2S U27790 ( .I1(n26534), .I2(n26048), .O(n26049) );
  MUX2 U27791 ( .A(n26049), .B(img[1189]), .S(n29207), .O(n12343) );
  BUF12CK U27792 ( .I(n26583), .O(n26534) );
  AOI22S U27793 ( .A1(n28037), .A2(n30779), .B1(n26091), .B2(img[1189]), .O(
        n26051) );
  ND2S U27794 ( .I1(n13820), .I2(img[1253]), .O(n26050) );
  ND3S U27795 ( .I1(n26534), .I2(n26051), .I3(n26050), .O(n26052) );
  MUX2 U27796 ( .A(img[1245]), .B(n26052), .S(n29211), .O(n12289) );
  AOI22S U27797 ( .A1(n28382), .A2(img[1253]), .B1(n23941), .B2(n30780), .O(
        n26053) );
  ND2S U27798 ( .I1(n26534), .I2(n26053), .O(n26054) );
  MUX2 U27799 ( .A(img[1181]), .B(n26054), .S(n29214), .O(n12353) );
  AOI22S U27800 ( .A1(n29407), .A2(n30781), .B1(n26091), .B2(img[1181]), .O(
        n26056) );
  ND3S U27801 ( .I1(n26534), .I2(n26056), .I3(n26055), .O(n26057) );
  MUX2 U27802 ( .A(img[1253]), .B(n26057), .S(n29218), .O(n12279) );
  AOI22S U27803 ( .A1(n28382), .A2(img[1373]), .B1(n13779), .B2(n30782), .O(
        n26058) );
  ND2S U27804 ( .I1(n26534), .I2(n26058), .O(n26059) );
  MUX2 U27805 ( .A(n26059), .B(img[1317]), .S(n29233), .O(n12217) );
  AOI22S U27806 ( .A1(n28075), .A2(n30783), .B1(n26091), .B2(img[1317]), .O(
        n26061) );
  ND3S U27807 ( .I1(n26534), .I2(n26061), .I3(n26060), .O(n26062) );
  MUX2 U27808 ( .A(img[1373]), .B(n26062), .S(n29237), .O(n12159) );
  AOI22S U27809 ( .A1(n28382), .A2(img[1381]), .B1(n24193), .B2(n30784), .O(
        n26063) );
  ND2S U27810 ( .I1(n26534), .I2(n26063), .O(n26064) );
  MUX2 U27811 ( .A(img[1309]), .B(n26064), .S(n29240), .O(n12223) );
  AOI22S U27812 ( .A1(n25062), .A2(n30785), .B1(n26091), .B2(img[1309]), .O(
        n26066) );
  ND3S U27813 ( .I1(n26534), .I2(n26066), .I3(n26065), .O(n26067) );
  MUX2 U27814 ( .A(img[1381]), .B(n26067), .S(n29245), .O(n12153) );
  AOI22S U27815 ( .A1(n28382), .A2(img[997]), .B1(n24193), .B2(n30786), .O(
        n26068) );
  ND2S U27816 ( .I1(n26534), .I2(n26068), .O(n26069) );
  MUX2 U27817 ( .A(img[925]), .B(n26069), .S(n29221), .O(n12609) );
  AOI22S U27818 ( .A1(n28382), .A2(img[925]), .B1(n28433), .B2(n30787), .O(
        n26070) );
  ND2S U27819 ( .I1(n26534), .I2(n26070), .O(n26071) );
  MUX2 U27820 ( .A(img[997]), .B(n26071), .S(n29224), .O(n12535) );
  AOI22S U27821 ( .A1(n28083), .A2(img[229]), .B1(n23918), .B2(n30788), .O(
        n26072) );
  ND2S U27822 ( .I1(n26534), .I2(n26072), .O(n26073) );
  MUX2 U27823 ( .A(img[157]), .B(n26073), .S(n29264), .O(n13377) );
  AOI22S U27824 ( .A1(n28083), .A2(img[157]), .B1(n25859), .B2(n30789), .O(
        n26074) );
  ND2S U27825 ( .I1(n26534), .I2(n26074), .O(n26075) );
  MUX2 U27826 ( .A(img[229]), .B(n26075), .S(n29267), .O(n13303) );
  AOI22S U27827 ( .A1(n28083), .A2(img[357]), .B1(n24374), .B2(n30790), .O(
        n26076) );
  ND2S U27828 ( .I1(n26534), .I2(n26076), .O(n26077) );
  AOI22S U27829 ( .A1(n28083), .A2(img[285]), .B1(n28182), .B2(n30791), .O(
        n26078) );
  ND2S U27830 ( .I1(n26534), .I2(n26078), .O(n26079) );
  MUX2 U27831 ( .A(img[357]), .B(n26079), .S(n29182), .O(n13177) );
  AOI22S U27832 ( .A1(n26101), .A2(img[485]), .B1(n28433), .B2(n30792), .O(
        n26080) );
  ND2S U27833 ( .I1(n26534), .I2(n26080), .O(n26081) );
  MUX2 U27834 ( .A(img[413]), .B(n26081), .S(n29270), .O(n13121) );
  AOI22S U27835 ( .A1(n26101), .A2(img[413]), .B1(n25591), .B2(n30793), .O(
        n26082) );
  ND2S U27836 ( .I1(n26534), .I2(n26082), .O(n26083) );
  MUX2 U27837 ( .A(img[485]), .B(n26083), .S(n29273), .O(n13047) );
  AOI22S U27838 ( .A1(n26101), .A2(img[1501]), .B1(n25377), .B2(n30794), .O(
        n26084) );
  ND2S U27839 ( .I1(n26534), .I2(n26084), .O(n26085) );
  MUX2 U27840 ( .A(n26085), .B(img[1445]), .S(n29248), .O(n12087) );
  AOI22S U27841 ( .A1(n28614), .A2(n30795), .B1(n26091), .B2(img[1445]), .O(
        n26087) );
  ND2S U27842 ( .I1(n13770), .I2(img[1509]), .O(n26086) );
  ND3S U27843 ( .I1(n26534), .I2(n26087), .I3(n26086), .O(n26088) );
  AOI22S U27844 ( .A1(n26101), .A2(img[1509]), .B1(n25859), .B2(n30796), .O(
        n26089) );
  ND2S U27845 ( .I1(n13807), .I2(n26089), .O(n26090) );
  MUX2 U27846 ( .A(n26090), .B(img[1437]), .S(n29255), .O(n12097) );
  AOI22S U27847 ( .A1(n28135), .A2(n26092), .B1(n26091), .B2(img[1437]), .O(
        n26094) );
  ND2S U27848 ( .I1(n13770), .I2(img[1501]), .O(n26093) );
  ND3S U27849 ( .I1(n26534), .I2(n26094), .I3(n26093), .O(n26095) );
  MUX2 U27850 ( .A(img[1509]), .B(n26095), .S(n29261), .O(n12023) );
  AOI22S U27851 ( .A1(n26101), .A2(img[869]), .B1(n28162), .B2(n30797), .O(
        n26096) );
  ND2S U27852 ( .I1(n26534), .I2(n26096), .O(n26097) );
  MUX2 U27853 ( .A(img[797]), .B(n26097), .S(n29227), .O(n12735) );
  INV1S U27854 ( .I(img[869]), .O(n26098) );
  AOI22S U27855 ( .A1(n26101), .A2(img[797]), .B1(n29242), .B2(n26098), .O(
        n26099) );
  ND2S U27856 ( .I1(n26534), .I2(n26099), .O(n26100) );
  MUX2 U27857 ( .A(n26100), .B(img[869]), .S(n29230), .O(n12665) );
  AOI22S U27858 ( .A1(n26101), .A2(img[741]), .B1(n28614), .B2(n30798), .O(
        n26102) );
  ND2S U27859 ( .I1(n26534), .I2(n26102), .O(n26103) );
  MUX2 U27860 ( .A(img[669]), .B(n26103), .S(n29201), .O(n12865) );
  AOI22S U27861 ( .A1(n25810), .A2(img[669]), .B1(n29096), .B2(n30799), .O(
        n26104) );
  ND2S U27862 ( .I1(n26534), .I2(n26104), .O(n26105) );
  AOI22S U27863 ( .A1(n28840), .A2(img[1861]), .B1(n28592), .B2(n30800), .O(
        n26106) );
  ND2S U27864 ( .I1(n26534), .I2(n26106), .O(n26107) );
  MUX2 U27865 ( .A(img[1853]), .B(n26107), .S(n28919), .O(n11679) );
  INV1S U27866 ( .I(img[1861]), .O(n26108) );
  AOI22S U27867 ( .A1(n28182), .A2(n26108), .B1(n24313), .B2(img[1853]), .O(
        n26110) );
  ND3S U27868 ( .I1(n26534), .I2(n26110), .I3(n26109), .O(n26111) );
  MUX2 U27869 ( .A(img[1861]), .B(n26111), .S(n28916), .O(n11673) );
  AOI22S U27870 ( .A1(n28106), .A2(img[1917]), .B1(n28182), .B2(n30801), .O(
        n26112) );
  ND2S U27871 ( .I1(n26534), .I2(n26112), .O(n26113) );
  AOI22S U27872 ( .A1(n28182), .A2(n30802), .B1(n28069), .B2(img[1797]), .O(
        n26115) );
  AOI22S U27873 ( .A1(n13905), .A2(img[1861]), .B1(img[1893]), .B2(n28908), 
        .O(n26114) );
  ND3S U27874 ( .I1(n26534), .I2(n26115), .I3(n26114), .O(n26116) );
  MUX2 U27875 ( .A(img[1917]), .B(n26116), .S(n28911), .O(n11615) );
  AOI22S U27876 ( .A1(n26970), .A2(img[1885]), .B1(n28343), .B2(n30803), .O(
        n26117) );
  ND2S U27877 ( .I1(n26534), .I2(n26117), .O(n26118) );
  INV1S U27878 ( .I(img[1885]), .O(n26119) );
  AOI22S U27879 ( .A1(n28182), .A2(n26119), .B1(n28069), .B2(img[1829]), .O(
        n26121) );
  ND2S U27880 ( .I1(n29124), .I2(img[1893]), .O(n26120) );
  ND3S U27881 ( .I1(n26534), .I2(n26121), .I3(n26120), .O(n26122) );
  MUX2 U27882 ( .A(img[1885]), .B(n26122), .S(n28896), .O(n11647) );
  AOI22S U27883 ( .A1(n28083), .A2(img[1893]), .B1(n27511), .B2(n30804), .O(
        n26123) );
  ND2S U27884 ( .I1(n26534), .I2(n26123), .O(n26124) );
  MUX2 U27885 ( .A(img[1821]), .B(n26124), .S(n28899), .O(n11711) );
  AOI22S U27886 ( .A1(n25062), .A2(n30805), .B1(n24313), .B2(img[1821]), .O(
        n26126) );
  AOI22S U27887 ( .A1(n13904), .A2(img[1885]), .B1(img[1917]), .B2(n13782), 
        .O(n26125) );
  ND3S U27888 ( .I1(n26534), .I2(n26126), .I3(n26125), .O(n26127) );
  MUX2 U27889 ( .A(img[1893]), .B(n26127), .S(n28903), .O(n11641) );
  AOI22S U27890 ( .A1(n28083), .A2(img[1733]), .B1(n25062), .B2(n30806), .O(
        n26128) );
  ND2S U27891 ( .I1(n26534), .I2(n26128), .O(n26129) );
  AOI22S U27892 ( .A1(n28592), .A2(n30807), .B1(n24313), .B2(img[1725]), .O(
        n26131) );
  ND2S U27893 ( .I1(n13770), .I2(img[1789]), .O(n26130) );
  ND3S U27894 ( .I1(n26534), .I2(n26131), .I3(n26130), .O(n26132) );
  MUX2 U27895 ( .A(img[1733]), .B(n26132), .S(n28945), .O(n11799) );
  AOI22S U27896 ( .A1(n28083), .A2(img[1789]), .B1(n25062), .B2(n30808), .O(
        n26133) );
  ND2S U27897 ( .I1(n26534), .I2(n26133), .O(n26134) );
  AOI22S U27898 ( .A1(n25377), .A2(n30809), .B1(n28069), .B2(img[1669]), .O(
        n26136) );
  AOI22S U27899 ( .A1(n13904), .A2(img[1733]), .B1(img[1765]), .B2(n13782), 
        .O(n26135) );
  ND3 U27900 ( .I1(n26583), .I2(n26136), .I3(n26135), .O(n26137) );
  AOI22S U27901 ( .A1(n28083), .A2(img[1757]), .B1(n28343), .B2(n30810), .O(
        n26138) );
  ND2S U27902 ( .I1(n26534), .I2(n26138), .O(n26139) );
  MUX2 U27903 ( .A(n26139), .B(img[1701]), .S(n28922), .O(n11831) );
  AOI22S U27904 ( .A1(n28862), .A2(n30811), .B1(n28043), .B2(img[1701]), .O(
        n26141) );
  ND2S U27905 ( .I1(n13770), .I2(img[1765]), .O(n26140) );
  ND3S U27906 ( .I1(n26534), .I2(n26141), .I3(n26140), .O(n26142) );
  AOI22S U27907 ( .A1(n28083), .A2(img[1765]), .B1(n13781), .B2(n30812), .O(
        n26143) );
  ND2S U27908 ( .I1(n26534), .I2(n26143), .O(n26144) );
  MUX2 U27909 ( .A(img[1693]), .B(n26144), .S(n28929), .O(n11841) );
  AOI22S U27910 ( .A1(n27735), .A2(n30813), .B1(n28069), .B2(img[1693]), .O(
        n26146) );
  AOI22S U27911 ( .A1(n13905), .A2(img[1757]), .B1(img[1789]), .B2(n13782), 
        .O(n26145) );
  ND3S U27912 ( .I1(n26534), .I2(n26146), .I3(n26145), .O(n26147) );
  MUX2 U27913 ( .A(img[1765]), .B(n26147), .S(n28933), .O(n11767) );
  AOI22S U27914 ( .A1(n28083), .A2(img[1605]), .B1(n28862), .B2(n30814), .O(
        n26148) );
  ND2S U27915 ( .I1(n26534), .I2(n26148), .O(n26149) );
  AOI22S U27916 ( .A1(n28075), .A2(n26150), .B1(n28069), .B2(img[1597]), .O(
        n26152) );
  ND2S U27917 ( .I1(n13770), .I2(img[1661]), .O(n26151) );
  ND3S U27918 ( .I1(n26534), .I2(n26152), .I3(n26151), .O(n26153) );
  MUX2 U27919 ( .A(img[1605]), .B(n26153), .S(n28973), .O(n11929) );
  AOI22S U27920 ( .A1(n28083), .A2(img[1661]), .B1(n27511), .B2(n30815), .O(
        n26154) );
  ND2S U27921 ( .I1(n26534), .I2(n26154), .O(n26155) );
  AOI22S U27922 ( .A1(n28075), .A2(n30816), .B1(n28069), .B2(img[1541]), .O(
        n26157) );
  AOI22S U27923 ( .A1(n13770), .A2(img[1605]), .B1(img[1637]), .B2(n13782), 
        .O(n26156) );
  ND3S U27924 ( .I1(n26534), .I2(n26157), .I3(n26156), .O(n26158) );
  MUX2 U27925 ( .A(img[1661]), .B(n26158), .S(n28969), .O(n11871) );
  AOI22S U27926 ( .A1(n28347), .A2(img[1629]), .B1(n27511), .B2(n30817), .O(
        n26159) );
  ND2S U27927 ( .I1(n26534), .I2(n26159), .O(n26160) );
  MUX2 U27928 ( .A(n26160), .B(img[1573]), .S(n28951), .O(n11961) );
  AOI22S U27929 ( .A1(n28592), .A2(n30818), .B1(n24313), .B2(img[1573]), .O(
        n26162) );
  ND3S U27930 ( .I1(n26534), .I2(n26162), .I3(n26161), .O(n26163) );
  AOI22S U27931 ( .A1(n26970), .A2(img[1637]), .B1(n13781), .B2(n30819), .O(
        n26164) );
  ND2S U27932 ( .I1(n26534), .I2(n26164), .O(n26165) );
  MUX2 U27933 ( .A(img[1565]), .B(n26165), .S(n28958), .O(n11967) );
  AOI22S U27934 ( .A1(n28037), .A2(n26166), .B1(n27919), .B2(img[1565]), .O(
        n26168) );
  AOI22S U27935 ( .A1(n13903), .A2(img[1629]), .B1(img[1661]), .B2(n13782), 
        .O(n26167) );
  ND3S U27936 ( .I1(n26534), .I2(n26168), .I3(n26167), .O(n26169) );
  MUX2 U27937 ( .A(img[1637]), .B(n26169), .S(n28962), .O(n11896) );
  AOI22S U27938 ( .A1(n28083), .A2(img[1117]), .B1(n27511), .B2(n30820), .O(
        n26170) );
  ND2S U27939 ( .I1(n26534), .I2(n26170), .O(n26171) );
  MUX2 U27940 ( .A(n26171), .B(img[1061]), .S(n29185), .O(n12473) );
  AOI22S U27941 ( .A1(n13781), .A2(n30821), .B1(n24946), .B2(img[1061]), .O(
        n26173) );
  ND3S U27942 ( .I1(n26534), .I2(n26173), .I3(n26172), .O(n26174) );
  MUX2 U27943 ( .A(img[1117]), .B(n26174), .S(n29189), .O(n12415) );
  AOI22S U27944 ( .A1(n25810), .A2(img[1125]), .B1(n27511), .B2(n30822), .O(
        n26175) );
  ND2S U27945 ( .I1(n26534), .I2(n26175), .O(n26176) );
  AOI22S U27946 ( .A1(n28075), .A2(n30823), .B1(n25444), .B2(img[1053]), .O(
        n26178) );
  ND3S U27947 ( .I1(n26534), .I2(n26178), .I3(n26177), .O(n26179) );
  MUX2 U27948 ( .A(img[1125]), .B(n26179), .S(n29198), .O(n12409) );
  AOI22S U27949 ( .A1(n28347), .A2(img[1989]), .B1(n29530), .B2(n30824), .O(
        n26180) );
  ND2S U27950 ( .I1(n26534), .I2(n26180), .O(n26181) );
  MUX2 U27951 ( .A(img[1981]), .B(n26181), .S(n29018), .O(n11553) );
  AOI22S U27952 ( .A1(n29242), .A2(n30825), .B1(n24434), .B2(img[1981]), .O(
        n26183) );
  ND2S U27953 ( .I1(n13770), .I2(img[2045]), .O(n26182) );
  ND3S U27954 ( .I1(n26534), .I2(n26183), .I3(n26182), .O(n26184) );
  MUX2 U27955 ( .A(img[1989]), .B(n26184), .S(n29015), .O(n11543) );
  AOI22S U27956 ( .A1(n28106), .A2(img[2045]), .B1(n24755), .B2(n30826), .O(
        n26185) );
  ND2S U27957 ( .I1(n26534), .I2(n26185), .O(n26186) );
  AOI22S U27958 ( .A1(n28135), .A2(n30827), .B1(n24313), .B2(img[1925]), .O(
        n26188) );
  AOI22S U27959 ( .A1(n29124), .A2(img[1989]), .B1(img[2021]), .B2(n13782), 
        .O(n26187) );
  ND3S U27960 ( .I1(n26534), .I2(n26188), .I3(n26187), .O(n26189) );
  MUX2 U27961 ( .A(img[2045]), .B(n26189), .S(n29011), .O(n11487) );
  AOI22S U27962 ( .A1(n25810), .A2(img[2013]), .B1(n24193), .B2(n30828), .O(
        n26190) );
  ND2S U27963 ( .I1(n26534), .I2(n26190), .O(n26191) );
  MUX2 U27964 ( .A(n26191), .B(img[1957]), .S(n28993), .O(n11575) );
  AOI22S U27965 ( .A1(n28135), .A2(n30829), .B1(n27919), .B2(img[1957]), .O(
        n26193) );
  ND3S U27966 ( .I1(n26534), .I2(n26193), .I3(n26192), .O(n26194) );
  AOI22S U27967 ( .A1(n24415), .A2(img[2021]), .B1(n28862), .B2(n30830), .O(
        n26195) );
  ND2S U27968 ( .I1(n26534), .I2(n26195), .O(n26196) );
  MUX2 U27969 ( .A(img[1949]), .B(n26196), .S(n29000), .O(n11585) );
  AOI22S U27970 ( .A1(n28135), .A2(n30831), .B1(n24946), .B2(img[1949]), .O(
        n26198) );
  AOI22S U27971 ( .A1(n29258), .A2(img[2013]), .B1(img[2045]), .B2(n28908), 
        .O(n26197) );
  ND3S U27972 ( .I1(n26534), .I2(n26198), .I3(n26197), .O(n26199) );
  MUX2 U27973 ( .A(img[2021]), .B(n26199), .S(n29004), .O(n11511) );
  AOI22S U27974 ( .A1(n27990), .A2(img[533]), .B1(n23918), .B2(n30832), .O(
        n26200) );
  ND2S U27975 ( .I1(n26534), .I2(n26200), .O(n26201) );
  MUX2 U27976 ( .A(n26201), .B(img[621]), .S(n29024), .O(n12911) );
  AOI22S U27977 ( .A1(n13776), .A2(img[621]), .B1(n23941), .B2(n30833), .O(
        n26202) );
  ND2S U27978 ( .I1(n26534), .I2(n26202), .O(n26203) );
  AOI22S U27979 ( .A1(n28442), .A2(img[21]), .B1(n24193), .B2(n30834), .O(
        n26204) );
  ND2S U27980 ( .I1(n26534), .I2(n26204), .O(n26205) );
  MUX2 U27981 ( .A(img[109]), .B(n26205), .S(n29030), .O(n13423) );
  AOI22S U27982 ( .A1(n13778), .A2(img[109]), .B1(n23941), .B2(n30835), .O(
        n26206) );
  ND2S U27983 ( .I1(n26534), .I2(n26206), .O(n26207) );
  AOI22S U27984 ( .A1(n13778), .A2(img[1237]), .B1(n28938), .B2(n30836), .O(
        n26208) );
  ND2S U27985 ( .I1(n26534), .I2(n26208), .O(n26209) );
  MUX2 U27986 ( .A(img[1197]), .B(n26209), .S(n29033), .O(n12337) );
  AOI22S U27987 ( .A1(n28135), .A2(n30837), .B1(n24313), .B2(img[1197]), .O(
        n26211) );
  ND3S U27988 ( .I1(n26534), .I2(n26211), .I3(n26210), .O(n26212) );
  MUX2 U27989 ( .A(img[1237]), .B(n26212), .S(n29037), .O(n12295) );
  AOI22S U27990 ( .A1(n13781), .A2(n30838), .B1(n24946), .B2(img[1173]), .O(
        n26214) );
  ND2S U27991 ( .I1(n13903), .I2(img[1237]), .O(n26213) );
  ND3S U27992 ( .I1(n26534), .I2(n26214), .I3(n26213), .O(n26215) );
  MUX2 U27993 ( .A(img[1261]), .B(n26215), .S(n29044), .O(n12273) );
  AOI22S U27994 ( .A1(n13778), .A2(img[1261]), .B1(n25062), .B2(n30839), .O(
        n26216) );
  ND2S U27995 ( .I1(n26534), .I2(n26216), .O(n26217) );
  AOI22S U27996 ( .A1(n13778), .A2(img[1365]), .B1(n28862), .B2(n30840), .O(
        n26218) );
  ND2S U27997 ( .I1(n26534), .I2(n26218), .O(n26219) );
  AOI22S U27998 ( .A1(n28162), .A2(n30841), .B1(n25444), .B2(img[1325]), .O(
        n26221) );
  ND2S U27999 ( .I1(n13770), .I2(img[1389]), .O(n26220) );
  ND3S U28000 ( .I1(n26534), .I2(n26221), .I3(n26220), .O(n26222) );
  MUX2 U28001 ( .A(img[1365]), .B(n26222), .S(n29051), .O(n12169) );
  AOI22S U28002 ( .A1(n28162), .A2(n30842), .B1(n24946), .B2(img[1301]), .O(
        n26224) );
  ND2S U28003 ( .I1(n13770), .I2(img[1365]), .O(n26223) );
  ND3S U28004 ( .I1(n26534), .I2(n26224), .I3(n26223), .O(n26225) );
  MUX2 U28005 ( .A(img[1389]), .B(n26225), .S(n29058), .O(n12143) );
  AOI22S U28006 ( .A1(n25595), .A2(img[1389]), .B1(n25377), .B2(n30843), .O(
        n26226) );
  ND2S U28007 ( .I1(n26534), .I2(n26226), .O(n26227) );
  MUX2 U28008 ( .A(n26227), .B(img[1301]), .S(n29054), .O(n12233) );
  AOI22S U28009 ( .A1(n24415), .A2(img[917]), .B1(n29096), .B2(n30844), .O(
        n26228) );
  ND2S U28010 ( .I1(n26534), .I2(n26228), .O(n26229) );
  MUX2 U28011 ( .A(img[1005]), .B(n26229), .S(n29064), .O(n12529) );
  AOI22S U28012 ( .A1(n28106), .A2(img[1005]), .B1(n28938), .B2(n30845), .O(
        n26230) );
  ND2S U28013 ( .I1(n26534), .I2(n26230), .O(n26231) );
  AOI22S U28014 ( .A1(n29072), .A2(img[149]), .B1(n29096), .B2(n30846), .O(
        n26232) );
  ND2S U28015 ( .I1(n26534), .I2(n26232), .O(n26233) );
  MUX2 U28016 ( .A(img[237]), .B(n26233), .S(n29070), .O(n13297) );
  AOI22S U28017 ( .A1(n13771), .A2(img[237]), .B1(n25377), .B2(n30847), .O(
        n26234) );
  ND2S U28018 ( .I1(n26534), .I2(n26234), .O(n26235) );
  MUX2 U28019 ( .A(img[149]), .B(n26235), .S(n29067), .O(n13383) );
  AOI22S U28020 ( .A1(n28106), .A2(img[277]), .B1(n25591), .B2(n30848), .O(
        n26236) );
  ND2S U28021 ( .I1(n26534), .I2(n26236), .O(n26237) );
  MUX2 U28022 ( .A(img[365]), .B(n26237), .S(n29078), .O(n13167) );
  AOI22S U28023 ( .A1(n24415), .A2(img[365]), .B1(n25062), .B2(n30849), .O(
        n26238) );
  ND2S U28024 ( .I1(n13807), .I2(n26238), .O(n26239) );
  AOI22S U28025 ( .A1(n13771), .A2(img[405]), .B1(n29096), .B2(n30850), .O(
        n26240) );
  ND2S U28026 ( .I1(n13807), .I2(n26240), .O(n26241) );
  MUX2 U28027 ( .A(img[493]), .B(n26241), .S(n29084), .O(n13041) );
  AOI22S U28028 ( .A1(n13780), .A2(img[493]), .B1(n25377), .B2(n30851), .O(
        n26242) );
  ND2S U28029 ( .I1(n13807), .I2(n26242), .O(n26243) );
  AOI22S U28030 ( .A1(n13780), .A2(img[1493]), .B1(n13781), .B2(n30852), .O(
        n26244) );
  ND2S U28031 ( .I1(n13807), .I2(n26244), .O(n26245) );
  AOI22S U28032 ( .A1(n25377), .A2(n30853), .B1(n24313), .B2(img[1453]), .O(
        n26247) );
  ND2S U28033 ( .I1(n13770), .I2(img[1517]), .O(n26246) );
  ND3S U28034 ( .I1(n26534), .I2(n26247), .I3(n26246), .O(n26248) );
  MUX2 U28035 ( .A(n26248), .B(img[1493]), .S(n29091), .O(n12039) );
  AOI22S U28036 ( .A1(n23941), .A2(n30854), .B1(n24313), .B2(img[1429]), .O(
        n26250) );
  ND2S U28037 ( .I1(n13770), .I2(img[1493]), .O(n26249) );
  ND3S U28038 ( .I1(n26534), .I2(n26250), .I3(n26249), .O(n26251) );
  AOI22S U28039 ( .A1(n13776), .A2(img[1517]), .B1(n28037), .B2(n30855), .O(
        n26252) );
  ND2S U28040 ( .I1(n13807), .I2(n26252), .O(n26253) );
  MUX2 U28041 ( .A(img[1429]), .B(n26253), .S(n29094), .O(n12103) );
  INV1S U28042 ( .I(img[877]), .O(n26254) );
  AOI22S U28043 ( .A1(n13778), .A2(img[789]), .B1(n29096), .B2(n26254), .O(
        n26255) );
  ND2S U28044 ( .I1(n13807), .I2(n26255), .O(n26256) );
  MUX2 U28045 ( .A(n26256), .B(img[877]), .S(n29106), .O(n12655) );
  AOI22S U28046 ( .A1(n13778), .A2(img[877]), .B1(n29194), .B2(n30856), .O(
        n26257) );
  ND2S U28047 ( .I1(n13807), .I2(n26257), .O(n26258) );
  AOI22S U28048 ( .A1(n13778), .A2(img[661]), .B1(n29096), .B2(n30857), .O(
        n26259) );
  ND2S U28049 ( .I1(n13807), .I2(n26259), .O(n26260) );
  MUX2 U28050 ( .A(n26260), .B(img[749]), .S(n29112), .O(n12785) );
  AOI22S U28051 ( .A1(n13778), .A2(img[749]), .B1(n25377), .B2(n30858), .O(
        n26261) );
  ND2S U28052 ( .I1(n13807), .I2(n26261), .O(n26262) );
  AOI22S U28053 ( .A1(n13778), .A2(img[1869]), .B1(n23941), .B2(n30859), .O(
        n26263) );
  ND2S U28054 ( .I1(n13807), .I2(n26263), .O(n26264) );
  MUX2 U28055 ( .A(n26264), .B(img[1845]), .S(n28693), .O(n11689) );
  AOI22S U28056 ( .A1(n28162), .A2(n30860), .B1(n28069), .B2(img[1845]), .O(
        n26266) );
  ND3S U28057 ( .I1(n26534), .I2(n26266), .I3(n26265), .O(n26267) );
  MUX2 U28058 ( .A(img[1869]), .B(n26267), .S(n28698), .O(n11663) );
  AOI22S U28059 ( .A1(n13778), .A2(img[1909]), .B1(n28913), .B2(n30861), .O(
        n26268) );
  ND2S U28060 ( .I1(n13807), .I2(n26268), .O(n26269) );
  AOI22S U28061 ( .A1(n28037), .A2(n30862), .B1(n24890), .B2(img[1805]), .O(
        n26271) );
  AOI22S U28062 ( .A1(n13903), .A2(img[1869]), .B1(img[1901]), .B2(n13782), 
        .O(n26270) );
  ND3S U28063 ( .I1(n26534), .I2(n26271), .I3(n26270), .O(n26272) );
  MUX2 U28064 ( .A(img[1909]), .B(n26272), .S(n28690), .O(n11625) );
  AOI22S U28065 ( .A1(n13778), .A2(img[1877]), .B1(n29407), .B2(n30863), .O(
        n26273) );
  ND2S U28066 ( .I1(n13807), .I2(n26273), .O(n26274) );
  MUX2 U28067 ( .A(n26274), .B(img[1837]), .S(n28672), .O(n11695) );
  AOI22S U28068 ( .A1(n28037), .A2(n30864), .B1(n24313), .B2(img[1837]), .O(
        n26276) );
  ND3S U28069 ( .I1(n26534), .I2(n26276), .I3(n26275), .O(n26277) );
  MUX2 U28070 ( .A(img[1877]), .B(n26277), .S(n28676), .O(n11657) );
  AOI22S U28071 ( .A1(n28862), .A2(n30865), .B1(n28069), .B2(img[1813]), .O(
        n26279) );
  AOI22S U28072 ( .A1(n29258), .A2(img[1877]), .B1(img[1909]), .B2(n13782), 
        .O(n26278) );
  ND3S U28073 ( .I1(n26534), .I2(n26279), .I3(n26278), .O(n26280) );
  MUX2 U28074 ( .A(img[1901]), .B(n26280), .S(n28683), .O(n11631) );
  AOI22S U28075 ( .A1(n29435), .A2(img[1901]), .B1(n29407), .B2(n30866), .O(
        n26281) );
  ND2S U28076 ( .I1(n13807), .I2(n26281), .O(n26282) );
  MUX2 U28077 ( .A(n26282), .B(img[1813]), .S(n28679), .O(n11721) );
  AOI22S U28078 ( .A1(n29129), .A2(img[1741]), .B1(n29397), .B2(n30867), .O(
        n26283) );
  ND2S U28079 ( .I1(n13807), .I2(n26283), .O(n26284) );
  MUX2 U28080 ( .A(n26284), .B(img[1717]), .S(n28722), .O(n11815) );
  AOI22S U28081 ( .A1(n13779), .A2(n30868), .B1(n26091), .B2(img[1717]), .O(
        n26286) );
  ND3S U28082 ( .I1(n26534), .I2(n26286), .I3(n26285), .O(n26287) );
  MUX2 U28083 ( .A(img[1741]), .B(n26287), .S(n28726), .O(n11793) );
  AOI22S U28084 ( .A1(n26101), .A2(img[1781]), .B1(n28913), .B2(n30869), .O(
        n26288) );
  ND2S U28085 ( .I1(n13807), .I2(n26288), .O(n26289) );
  MUX2 U28086 ( .A(img[1677]), .B(n26289), .S(n28715), .O(n11857) );
  AOI22S U28087 ( .A1(n28343), .A2(n30870), .B1(n27919), .B2(img[1677]), .O(
        n26291) );
  AOI22S U28088 ( .A1(n13770), .A2(img[1741]), .B1(img[1773]), .B2(n28908), 
        .O(n26290) );
  ND3S U28089 ( .I1(n26534), .I2(n26291), .I3(n26290), .O(n26292) );
  MUX2 U28090 ( .A(img[1781]), .B(n26292), .S(n28719), .O(n11751) );
  AOI22S U28091 ( .A1(n13771), .A2(img[1749]), .B1(n25591), .B2(n30871), .O(
        n26293) );
  ND2S U28092 ( .I1(n13807), .I2(n26293), .O(n26294) );
  MUX2 U28093 ( .A(n26294), .B(img[1709]), .S(n28701), .O(n11825) );
  AOI22S U28094 ( .A1(n25591), .A2(n30872), .B1(n27919), .B2(img[1709]), .O(
        n26296) );
  ND3S U28095 ( .I1(n26534), .I2(n26296), .I3(n26295), .O(n26297) );
  MUX2 U28096 ( .A(img[1749]), .B(n26297), .S(n28705), .O(n11783) );
  AOI22S U28097 ( .A1(n28938), .A2(n30873), .B1(n24313), .B2(img[1685]), .O(
        n26299) );
  AOI22S U28098 ( .A1(n13904), .A2(img[1749]), .B1(img[1781]), .B2(n28908), 
        .O(n26298) );
  ND3S U28099 ( .I1(n26534), .I2(n26299), .I3(n26298), .O(n26300) );
  MUX2 U28100 ( .A(img[1773]), .B(n26300), .S(n28712), .O(n11761) );
  AOI22S U28101 ( .A1(n13776), .A2(img[1773]), .B1(n25591), .B2(n30874), .O(
        n26301) );
  ND2S U28102 ( .I1(n13807), .I2(n26301), .O(n26302) );
  MUX2 U28103 ( .A(n26302), .B(img[1685]), .S(n28708), .O(n11847) );
  AOI22S U28104 ( .A1(n13771), .A2(img[1613]), .B1(n27511), .B2(n30875), .O(
        n26303) );
  ND2S U28105 ( .I1(n13807), .I2(n26303), .O(n26304) );
  MUX2 U28106 ( .A(n26304), .B(img[1589]), .S(n28750), .O(n11945) );
  AOI22S U28107 ( .A1(n25062), .A2(n30876), .B1(n27919), .B2(img[1589]), .O(
        n26306) );
  ND3S U28108 ( .I1(n26534), .I2(n26306), .I3(n26305), .O(n26307) );
  MUX2 U28109 ( .A(img[1613]), .B(n26307), .S(n28754), .O(n11919) );
  AOI22S U28110 ( .A1(n13778), .A2(img[1653]), .B1(n27511), .B2(n30877), .O(
        n26308) );
  ND2S U28111 ( .I1(n13807), .I2(n26308), .O(n26309) );
  AOI22S U28112 ( .A1(n28938), .A2(n30878), .B1(n24313), .B2(img[1549]), .O(
        n26311) );
  AOI22S U28113 ( .A1(n29258), .A2(img[1613]), .B1(img[1645]), .B2(n13782), 
        .O(n26310) );
  ND3S U28114 ( .I1(n26534), .I2(n26311), .I3(n26310), .O(n26312) );
  MUX2 U28115 ( .A(img[1653]), .B(n26312), .S(n28747), .O(n11881) );
  AOI22S U28116 ( .A1(n13772), .A2(img[1621]), .B1(n27511), .B2(n30879), .O(
        n26313) );
  ND2S U28117 ( .I1(n13807), .I2(n26313), .O(n26314) );
  MUX2 U28118 ( .A(n26314), .B(img[1581]), .S(n28729), .O(n11951) );
  AOI22S U28119 ( .A1(n28938), .A2(n30880), .B1(n27919), .B2(img[1581]), .O(
        n26316) );
  ND3S U28120 ( .I1(n26534), .I2(n26316), .I3(n26315), .O(n26317) );
  MUX2 U28121 ( .A(img[1621]), .B(n26317), .S(n28733), .O(n11913) );
  AOI22S U28122 ( .A1(n28938), .A2(n30881), .B1(n27919), .B2(img[1557]), .O(
        n26319) );
  AOI22S U28123 ( .A1(n29258), .A2(img[1621]), .B1(img[1653]), .B2(n13782), 
        .O(n26318) );
  ND3S U28124 ( .I1(n26534), .I2(n26319), .I3(n26318), .O(n26320) );
  MUX2 U28125 ( .A(img[1645]), .B(n26320), .S(n28740), .O(n11887) );
  AOI22S U28126 ( .A1(n13780), .A2(img[1645]), .B1(n28037), .B2(n30882), .O(
        n26321) );
  ND2S U28127 ( .I1(n13807), .I2(n26321), .O(n26322) );
  MUX2 U28128 ( .A(n26322), .B(img[1557]), .S(n28736), .O(n11977) );
  AOI22S U28129 ( .A1(n13777), .A2(img[1109]), .B1(n27511), .B2(n30883), .O(
        n26323) );
  ND2S U28130 ( .I1(n13807), .I2(n26323), .O(n26324) );
  MUX2 U28131 ( .A(n26324), .B(img[1069]), .S(n29115), .O(n12463) );
  AOI22S U28132 ( .A1(n28938), .A2(n30884), .B1(n28254), .B2(img[1069]), .O(
        n26326) );
  ND2S U28133 ( .I1(n13902), .I2(img[1133]), .O(n26325) );
  ND3S U28134 ( .I1(n26534), .I2(n26326), .I3(n26325), .O(n26327) );
  MUX2 U28135 ( .A(img[1109]), .B(n26327), .S(n29119), .O(n12425) );
  AOI22S U28136 ( .A1(n28938), .A2(n30885), .B1(n28069), .B2(img[1045]), .O(
        n26329) );
  ND2S U28137 ( .I1(n13819), .I2(img[1109]), .O(n26328) );
  ND3S U28138 ( .I1(n26534), .I2(n26329), .I3(n26328), .O(n26330) );
  MUX2 U28139 ( .A(img[1133]), .B(n26330), .S(n29127), .O(n12399) );
  AOI22S U28140 ( .A1(n13778), .A2(img[1133]), .B1(n25859), .B2(n30886), .O(
        n26331) );
  ND2S U28141 ( .I1(n13807), .I2(n26331), .O(n26332) );
  MUX2 U28142 ( .A(n26332), .B(img[1045]), .S(n29122), .O(n12488) );
  AOI22S U28143 ( .A1(n25595), .A2(img[1997]), .B1(n13781), .B2(n30887), .O(
        n26333) );
  ND2S U28144 ( .I1(n13807), .I2(n26333), .O(n26334) );
  MUX2 U28145 ( .A(n26334), .B(img[1973]), .S(n28792), .O(n11559) );
  INV1S U28146 ( .I(img[1997]), .O(n26335) );
  AOI22S U28147 ( .A1(n28938), .A2(n26335), .B1(n24808), .B2(img[1973]), .O(
        n26337) );
  ND3S U28148 ( .I1(n26534), .I2(n26337), .I3(n26336), .O(n26338) );
  MUX2 U28149 ( .A(img[1997]), .B(n26338), .S(n28796), .O(n11537) );
  AOI22S U28150 ( .A1(n26101), .A2(img[2037]), .B1(n24755), .B2(n30888), .O(
        n26339) );
  ND2S U28151 ( .I1(n13807), .I2(n26339), .O(n26340) );
  MUX2 U28152 ( .A(img[1933]), .B(n26340), .S(n28785), .O(n11601) );
  AOI22S U28153 ( .A1(n25062), .A2(n30889), .B1(n27919), .B2(img[1933]), .O(
        n26342) );
  AOI22S U28154 ( .A1(n29258), .A2(img[1997]), .B1(img[2029]), .B2(n13782), 
        .O(n26341) );
  ND3S U28155 ( .I1(n26534), .I2(n26342), .I3(n26341), .O(n26343) );
  MUX2 U28156 ( .A(img[2037]), .B(n26343), .S(n28789), .O(n11495) );
  AOI22S U28157 ( .A1(n25810), .A2(img[2005]), .B1(n28433), .B2(n30890), .O(
        n26344) );
  ND2S U28158 ( .I1(n13807), .I2(n26344), .O(n26345) );
  AOI22S U28159 ( .A1(n25591), .A2(n30891), .B1(n28069), .B2(img[1965]), .O(
        n26347) );
  ND2S U28160 ( .I1(n29124), .I2(img[2029]), .O(n26346) );
  ND3S U28161 ( .I1(n26534), .I2(n26347), .I3(n26346), .O(n26348) );
  MUX2 U28162 ( .A(img[2005]), .B(n26348), .S(n28775), .O(n11527) );
  AOI22S U28163 ( .A1(n29194), .A2(n30892), .B1(n24313), .B2(img[1941]), .O(
        n26350) );
  AOI22S U28164 ( .A1(n13820), .A2(img[2005]), .B1(img[2037]), .B2(n13782), 
        .O(n26349) );
  ND3S U28165 ( .I1(n26534), .I2(n26350), .I3(n26349), .O(n26351) );
  MUX2 U28166 ( .A(img[2029]), .B(n26351), .S(n28782), .O(n11505) );
  AOI22S U28167 ( .A1(n26822), .A2(img[2029]), .B1(n23918), .B2(n30893), .O(
        n26352) );
  ND2S U28168 ( .I1(n13807), .I2(n26352), .O(n26353) );
  MUX2 U28169 ( .A(n26353), .B(img[1941]), .S(n28778), .O(n11591) );
  AOI22S U28170 ( .A1(n28347), .A2(img[197]), .B1(n24374), .B2(n30894), .O(
        n26354) );
  ND2S U28171 ( .I1(n13807), .I2(n26354), .O(n26355) );
  MUX2 U28172 ( .A(img[189]), .B(n26355), .S(n28848), .O(n13345) );
  AOI22S U28173 ( .A1(n28442), .A2(img[189]), .B1(n29096), .B2(n30895), .O(
        n26356) );
  ND2S U28174 ( .I1(n13807), .I2(n26356), .O(n26357) );
  MUX2 U28175 ( .A(img[197]), .B(n26357), .S(n28845), .O(n13335) );
  AOI22S U28176 ( .A1(n28347), .A2(img[69]), .B1(n27049), .B2(n30896), .O(
        n26358) );
  ND2S U28177 ( .I1(n13807), .I2(n26358), .O(n26359) );
  MUX2 U28178 ( .A(img[61]), .B(n26359), .S(n28807), .O(n13471) );
  AOI22S U28179 ( .A1(n28106), .A2(img[61]), .B1(n27049), .B2(n30897), .O(
        n26360) );
  ND2S U28180 ( .I1(n13807), .I2(n26360), .O(n26361) );
  MUX2 U28181 ( .A(img[69]), .B(n26361), .S(n28804), .O(n13465) );
  AOI22S U28182 ( .A1(n26970), .A2(img[1277]), .B1(n27049), .B2(n30898), .O(
        n26362) );
  ND2S U28183 ( .I1(n13807), .I2(n26362), .O(n26363) );
  INV1S U28184 ( .I(img[1277]), .O(n26364) );
  AOI22S U28185 ( .A1(n25062), .A2(n26364), .B1(n28043), .B2(img[1157]), .O(
        n26366) );
  ND2S U28186 ( .I1(n13902), .I2(img[1221]), .O(n26365) );
  ND3S U28187 ( .I1(n26534), .I2(n26366), .I3(n26365), .O(n26367) );
  MUX2 U28188 ( .A(img[1277]), .B(n26367), .S(n28814), .O(n12257) );
  AOI22S U28189 ( .A1(n28347), .A2(img[1221]), .B1(n25591), .B2(n30899), .O(
        n26368) );
  ND2S U28190 ( .I1(n13807), .I2(n26368), .O(n26369) );
  MUX2 U28191 ( .A(img[1213]), .B(n26369), .S(n28821), .O(n12321) );
  INV1S U28192 ( .I(img[1221]), .O(n26370) );
  AOI22S U28193 ( .A1(n28343), .A2(n26370), .B1(n24313), .B2(img[1213]), .O(
        n26372) );
  ND2S U28194 ( .I1(n13770), .I2(img[1277]), .O(n26371) );
  ND3S U28195 ( .I1(n26534), .I2(n26372), .I3(n26371), .O(n26373) );
  MUX2 U28196 ( .A(img[1221]), .B(n26373), .S(n28818), .O(n12311) );
  AOI22S U28197 ( .A1(n29072), .A2(img[1405]), .B1(n29530), .B2(n30900), .O(
        n26374) );
  ND2S U28198 ( .I1(n13807), .I2(n26374), .O(n26375) );
  INV1S U28199 ( .I(img[1405]), .O(n26376) );
  AOI22S U28200 ( .A1(n25062), .A2(n26376), .B1(n26504), .B2(img[1285]), .O(
        n26378) );
  ND3S U28201 ( .I1(n26534), .I2(n26378), .I3(n26377), .O(n26379) );
  MUX2 U28202 ( .A(img[1405]), .B(n26379), .S(n28828), .O(n12127) );
  AOI22S U28203 ( .A1(n29129), .A2(img[1349]), .B1(n29096), .B2(n30901), .O(
        n26380) );
  ND2S U28204 ( .I1(n13807), .I2(n26380), .O(n26381) );
  MUX2 U28205 ( .A(img[1341]), .B(n26381), .S(n28835), .O(n12191) );
  INV1S U28206 ( .I(img[1349]), .O(n26382) );
  AOI22S U28207 ( .A1(n28182), .A2(n26382), .B1(n26504), .B2(img[1341]), .O(
        n26384) );
  ND3S U28208 ( .I1(n26534), .I2(n26384), .I3(n26383), .O(n26385) );
  MUX2 U28209 ( .A(img[1349]), .B(n26385), .S(n28832), .O(n12185) );
  AOI22S U28210 ( .A1(n13778), .A2(img[965]), .B1(n13781), .B2(n30902), .O(
        n26386) );
  ND2S U28211 ( .I1(n13807), .I2(n26386), .O(n26387) );
  AOI22S U28212 ( .A1(n27065), .A2(img[957]), .B1(n28135), .B2(n30903), .O(
        n26388) );
  ND2S U28213 ( .I1(n13807), .I2(n26388), .O(n26389) );
  MUX2 U28214 ( .A(img[965]), .B(n26389), .S(n28838), .O(n12567) );
  AOI22S U28215 ( .A1(n28221), .A2(img[325]), .B1(n25062), .B2(n30904), .O(
        n26390) );
  ND2S U28216 ( .I1(n13807), .I2(n26390), .O(n26391) );
  AOI22S U28217 ( .A1(n27685), .A2(img[317]), .B1(n28913), .B2(n30905), .O(
        n26392) );
  ND2S U28218 ( .I1(n13807), .I2(n26392), .O(n26393) );
  MUX2 U28219 ( .A(img[325]), .B(n26393), .S(n28851), .O(n13209) );
  AOI22S U28220 ( .A1(n24415), .A2(img[453]), .B1(n24193), .B2(n30906), .O(
        n26394) );
  ND2S U28221 ( .I1(n13807), .I2(n26394), .O(n26395) );
  MUX2 U28222 ( .A(img[445]), .B(n26395), .S(n28860), .O(n13090) );
  AOI22S U28223 ( .A1(n28840), .A2(img[445]), .B1(n28862), .B2(n30907), .O(
        n26396) );
  ND2S U28224 ( .I1(n13807), .I2(n26396), .O(n26397) );
  MUX2 U28225 ( .A(img[453]), .B(n26397), .S(n28857), .O(n13079) );
  AOI22S U28226 ( .A1(n26101), .A2(img[1533]), .B1(n28182), .B2(n30908), .O(
        n26398) );
  ND2S U28227 ( .I1(n13807), .I2(n26398), .O(n26399) );
  AOI22S U28228 ( .A1(n25062), .A2(n30909), .B1(n26504), .B2(img[1413]), .O(
        n26401) );
  ND2S U28229 ( .I1(n13819), .I2(img[1477]), .O(n26400) );
  ND3S U28230 ( .I1(n26534), .I2(n26401), .I3(n26400), .O(n26402) );
  MUX2 U28231 ( .A(img[1533]), .B(n26402), .S(n28868), .O(n12001) );
  AOI22S U28232 ( .A1(n13771), .A2(img[1477]), .B1(n28913), .B2(n30910), .O(
        n26403) );
  ND2S U28233 ( .I1(n13807), .I2(n26403), .O(n26404) );
  MUX2 U28234 ( .A(img[1469]), .B(n26404), .S(n28875), .O(n12065) );
  AOI22S U28235 ( .A1(n28343), .A2(n30911), .B1(n26504), .B2(img[1469]), .O(
        n26406) );
  ND3 U28236 ( .I1(n26583), .I2(n26406), .I3(n26405), .O(n26407) );
  AOI22S U28237 ( .A1(n26101), .A2(img[837]), .B1(n27735), .B2(n30912), .O(
        n26408) );
  ND2S U28238 ( .I1(n13807), .I2(n26408), .O(n26409) );
  INV1S U28239 ( .I(img[837]), .O(n26410) );
  AOI22S U28240 ( .A1(n24415), .A2(img[829]), .B1(n13781), .B2(n26410), .O(
        n26411) );
  ND2S U28241 ( .I1(n13807), .I2(n26411), .O(n26412) );
  MUX2 U28242 ( .A(n26412), .B(img[837]), .S(n28879), .O(n12697) );
  AOI22S U28243 ( .A1(n28347), .A2(img[1149]), .B1(n13781), .B2(n30913), .O(
        n26413) );
  ND2S U28244 ( .I1(n13807), .I2(n26413), .O(n26414) );
  MUX2 U28245 ( .A(img[1029]), .B(n26414), .S(n28979), .O(n12505) );
  AOI22S U28246 ( .A1(n28343), .A2(n30914), .B1(n26504), .B2(img[1029]), .O(
        n26416) );
  ND3S U28247 ( .I1(n26534), .I2(n26416), .I3(n26415), .O(n26417) );
  MUX2 U28248 ( .A(img[1149]), .B(n26417), .S(n28983), .O(n12383) );
  AOI22S U28249 ( .A1(n28347), .A2(img[1093]), .B1(n13781), .B2(n30915), .O(
        n26418) );
  ND2S U28250 ( .I1(n13807), .I2(n26418), .O(n26419) );
  AOI22S U28251 ( .A1(n28343), .A2(n30916), .B1(n26504), .B2(img[1085]), .O(
        n26421) );
  ND2S U28252 ( .I1(n13820), .I2(img[1149]), .O(n26420) );
  ND3S U28253 ( .I1(n26534), .I2(n26421), .I3(n26420), .O(n26422) );
  MUX2 U28254 ( .A(img[1093]), .B(n26422), .S(n28987), .O(n12438) );
  AOI22S U28255 ( .A1(n28347), .A2(img[581]), .B1(n29242), .B2(n30917), .O(
        n26423) );
  ND2S U28256 ( .I1(n26534), .I2(n26423), .O(n26424) );
  MUX2 U28257 ( .A(n26424), .B(img[573]), .S(n29532), .O(n12959) );
  AOI22S U28258 ( .A1(n13772), .A2(img[573]), .B1(n27511), .B2(n30918), .O(
        n26425) );
  ND2S U28259 ( .I1(n26534), .I2(n26425), .O(n26426) );
  MUX2 U28260 ( .A(n26426), .B(img[581]), .S(n28799), .O(n12953) );
  AOI22S U28261 ( .A1(n13776), .A2(img[709]), .B1(n13781), .B2(n30919), .O(
        n26427) );
  ND2S U28262 ( .I1(n26534), .I2(n26427), .O(n26428) );
  AOI22S U28263 ( .A1(n25810), .A2(img[701]), .B1(n13781), .B2(n30920), .O(
        n26429) );
  ND2S U28264 ( .I1(n26534), .I2(n26429), .O(n26430) );
  AOI22S U28265 ( .A1(n26855), .A2(img[597]), .B1(n23941), .B2(n30921), .O(
        n26431) );
  ND2S U28266 ( .I1(n26534), .I2(n26431), .O(n26432) );
  MUX2 U28267 ( .A(n26432), .B(img[557]), .S(n29439), .O(n12975) );
  AOI22S U28268 ( .A1(n28347), .A2(img[557]), .B1(n28862), .B2(n30922), .O(
        n26433) );
  ND2S U28269 ( .I1(n26534), .I2(n26433), .O(n26434) );
  MUX2 U28270 ( .A(n26434), .B(img[597]), .S(n29133), .O(n12937) );
  AOI22S U28271 ( .A1(n28412), .A2(img[85]), .B1(n13781), .B2(n30923), .O(
        n26435) );
  ND2S U28272 ( .I1(n26534), .I2(n26435), .O(n26436) );
  MUX2 U28273 ( .A(img[45]), .B(n26436), .S(n29136), .O(n13487) );
  AOI22S U28274 ( .A1(n28347), .A2(img[45]), .B1(n28343), .B2(n30924), .O(
        n26437) );
  ND2S U28275 ( .I1(n26534), .I2(n26437), .O(n26438) );
  MUX2 U28276 ( .A(img[85]), .B(n26438), .S(n29139), .O(n13449) );
  AOI22S U28277 ( .A1(n28106), .A2(img[981]), .B1(n24193), .B2(n30925), .O(
        n26439) );
  ND2S U28278 ( .I1(n26534), .I2(n26439), .O(n26440) );
  AOI22S U28279 ( .A1(n26490), .A2(img[941]), .B1(n23918), .B2(n30926), .O(
        n26441) );
  ND2S U28280 ( .I1(n26534), .I2(n26441), .O(n26442) );
  MUX2 U28281 ( .A(img[981]), .B(n26442), .S(n29145), .O(n12551) );
  AOI22S U28282 ( .A1(n26490), .A2(img[213]), .B1(n28862), .B2(n30927), .O(
        n26443) );
  ND2S U28283 ( .I1(n26534), .I2(n26443), .O(n26444) );
  MUX2 U28284 ( .A(img[173]), .B(n26444), .S(n29148), .O(n13361) );
  AOI22S U28285 ( .A1(n26490), .A2(img[173]), .B1(n28162), .B2(n30928), .O(
        n26445) );
  ND2S U28286 ( .I1(n26534), .I2(n26445), .O(n26446) );
  MUX2 U28287 ( .A(img[213]), .B(n26446), .S(n29151), .O(n13319) );
  AOI22S U28288 ( .A1(n26490), .A2(img[341]), .B1(n24374), .B2(n30929), .O(
        n26447) );
  ND2S U28289 ( .I1(n26534), .I2(n26447), .O(n26448) );
  MUX2 U28290 ( .A(img[301]), .B(n26448), .S(n29154), .O(n13231) );
  AOI22S U28291 ( .A1(n28347), .A2(img[301]), .B1(n25591), .B2(n30930), .O(
        n26449) );
  ND2S U28292 ( .I1(n26534), .I2(n26449), .O(n26450) );
  AOI22S U28293 ( .A1(n26855), .A2(img[469]), .B1(n25591), .B2(n30931), .O(
        n26451) );
  ND2S U28294 ( .I1(n26534), .I2(n26451), .O(n26452) );
  MUX2 U28295 ( .A(img[429]), .B(n26452), .S(n29160), .O(n13105) );
  AOI22S U28296 ( .A1(n28347), .A2(img[429]), .B1(n23941), .B2(n30932), .O(
        n26453) );
  ND2S U28297 ( .I1(n26534), .I2(n26453), .O(n26454) );
  MUX2 U28298 ( .A(img[469]), .B(n26454), .S(n29163), .O(n13063) );
  AOI22S U28299 ( .A1(n28347), .A2(img[853]), .B1(n28343), .B2(n30933), .O(
        n26455) );
  ND2S U28300 ( .I1(n26534), .I2(n26455), .O(n26456) );
  AOI22S U28301 ( .A1(n28347), .A2(img[813]), .B1(n28075), .B2(n30934), .O(
        n26457) );
  ND2S U28302 ( .I1(n26534), .I2(n26457), .O(n26458) );
  MUX2 U28303 ( .A(n26458), .B(img[853]), .S(n29170), .O(n12681) );
  AOI22S U28304 ( .A1(n28347), .A2(img[725]), .B1(n28037), .B2(n30935), .O(
        n26459) );
  ND2S U28305 ( .I1(n26534), .I2(n26459), .O(n26460) );
  AOI22S U28306 ( .A1(n28347), .A2(img[685]), .B1(n25062), .B2(n30936), .O(
        n26461) );
  ND2S U28307 ( .I1(n26534), .I2(n26461), .O(n26462) );
  AOI22S U28308 ( .A1(n28347), .A2(img[333]), .B1(n13781), .B2(n30937), .O(
        n26463) );
  ND2S U28309 ( .I1(n26534), .I2(n26463), .O(n26464) );
  AOI22S U28310 ( .A1(n28643), .A2(img[309]), .B1(n29457), .B2(n30938), .O(
        n26465) );
  ND2S U28311 ( .I1(n26534), .I2(n26465), .O(n26466) );
  MUX2 U28312 ( .A(img[333]), .B(n26466), .S(n28635), .O(n13199) );
  AOI22S U28313 ( .A1(n13777), .A2(img[1141]), .B1(n28162), .B2(n30939), .O(
        n26467) );
  ND2S U28314 ( .I1(n26534), .I2(n26467), .O(n26468) );
  MUX2 U28315 ( .A(img[1037]), .B(n26468), .S(n28757), .O(n12495) );
  AOI22S U28316 ( .A1(n29194), .A2(n30940), .B1(n26504), .B2(img[1037]), .O(
        n26470) );
  ND2S U28317 ( .I1(n13905), .I2(img[1101]), .O(n26469) );
  ND3S U28318 ( .I1(n26534), .I2(n26470), .I3(n26469), .O(n26471) );
  MUX2 U28319 ( .A(img[1141]), .B(n26471), .S(n28761), .O(n12393) );
  AOI22S U28320 ( .A1(n28840), .A2(img[1101]), .B1(n24755), .B2(n30941), .O(
        n26472) );
  ND2S U28321 ( .I1(n26534), .I2(n26472), .O(n26473) );
  MUX2 U28322 ( .A(n26473), .B(img[1077]), .S(n28764), .O(n12457) );
  AOI22S U28323 ( .A1(n29194), .A2(n26474), .B1(n26504), .B2(img[1077]), .O(
        n26476) );
  ND3S U28324 ( .I1(n26534), .I2(n26476), .I3(n26475), .O(n26477) );
  MUX2 U28325 ( .A(img[1101]), .B(n26477), .S(n28768), .O(n12431) );
  AOI22S U28326 ( .A1(n26490), .A2(img[717]), .B1(n24755), .B2(n30942), .O(
        n26478) );
  ND2S U28327 ( .I1(n26534), .I2(n26478), .O(n26479) );
  AOI22S U28328 ( .A1(n26490), .A2(img[693]), .B1(n29397), .B2(n30943), .O(
        n26480) );
  ND2S U28329 ( .I1(n26534), .I2(n26480), .O(n26481) );
  AOI22S U28330 ( .A1(n26490), .A2(img[589]), .B1(n28695), .B2(n30944), .O(
        n26482) );
  ND2S U28331 ( .I1(n26534), .I2(n26482), .O(n26483) );
  MUX2 U28332 ( .A(n26483), .B(img[565]), .S(n28578), .O(n12969) );
  AOI22S U28333 ( .A1(n26490), .A2(img[565]), .B1(n28938), .B2(n30945), .O(
        n26484) );
  ND2S U28334 ( .I1(n26534), .I2(n26484), .O(n26485) );
  MUX2 U28335 ( .A(n26485), .B(img[589]), .S(n28581), .O(n12943) );
  AOI22S U28336 ( .A1(n26490), .A2(img[77]), .B1(n28938), .B2(n30946), .O(
        n26486) );
  ND2S U28337 ( .I1(n26534), .I2(n26486), .O(n26487) );
  MUX2 U28338 ( .A(img[53]), .B(n26487), .S(n28584), .O(n13478) );
  AOI22S U28339 ( .A1(n26490), .A2(img[53]), .B1(n24193), .B2(n30947), .O(
        n26488) );
  ND2S U28340 ( .I1(n26534), .I2(n26488), .O(n26489) );
  AOI22S U28341 ( .A1(n26490), .A2(img[1269]), .B1(n27049), .B2(n30948), .O(
        n26491) );
  ND2S U28342 ( .I1(n26534), .I2(n26491), .O(n26492) );
  AOI22S U28343 ( .A1(n28135), .A2(n30949), .B1(n26504), .B2(img[1165]), .O(
        n26494) );
  ND2S U28344 ( .I1(n13902), .I2(img[1229]), .O(n26493) );
  ND3S U28345 ( .I1(n26534), .I2(n26494), .I3(n26493), .O(n26495) );
  MUX2 U28346 ( .A(img[1269]), .B(n26495), .S(n28595), .O(n12263) );
  AOI22S U28347 ( .A1(n28412), .A2(img[1229]), .B1(n28938), .B2(n30950), .O(
        n26496) );
  ND2S U28348 ( .I1(n26534), .I2(n26496), .O(n26497) );
  AOI22S U28349 ( .A1(n28135), .A2(n26498), .B1(n26504), .B2(img[1205]), .O(
        n26500) );
  ND2S U28350 ( .I1(n29124), .I2(img[1269]), .O(n26499) );
  ND3S U28351 ( .I1(n26534), .I2(n26500), .I3(n26499), .O(n26501) );
  MUX2 U28352 ( .A(img[1229]), .B(n26501), .S(n28602), .O(n12305) );
  AOI22S U28353 ( .A1(n28412), .A2(img[1397]), .B1(n28938), .B2(n30951), .O(
        n26502) );
  ND2S U28354 ( .I1(n26534), .I2(n26502), .O(n26503) );
  MUX2 U28355 ( .A(img[1293]), .B(n26503), .S(n28605), .O(n12239) );
  AOI22S U28356 ( .A1(n28075), .A2(n30952), .B1(n26504), .B2(img[1293]), .O(
        n26506) );
  ND3S U28357 ( .I1(n26534), .I2(n26506), .I3(n26505), .O(n26507) );
  MUX2 U28358 ( .A(img[1397]), .B(n26507), .S(n28609), .O(n12137) );
  AOI22S U28359 ( .A1(n25595), .A2(img[1357]), .B1(n25062), .B2(n30953), .O(
        n26508) );
  ND2S U28360 ( .I1(n26534), .I2(n26508), .O(n26509) );
  MUX2 U28361 ( .A(n26509), .B(img[1333]), .S(n28612), .O(n12201) );
  AOI22S U28362 ( .A1(n27443), .A2(n30954), .B1(n28069), .B2(img[1333]), .O(
        n26511) );
  ND2S U28363 ( .I1(n13819), .I2(img[1397]), .O(n26510) );
  ND3S U28364 ( .I1(n26534), .I2(n26511), .I3(n26510), .O(n26512) );
  MUX2 U28365 ( .A(img[1357]), .B(n26512), .S(n28617), .O(n12175) );
  AOI22S U28366 ( .A1(n28347), .A2(img[973]), .B1(n29194), .B2(n30955), .O(
        n26513) );
  ND2S U28367 ( .I1(n26534), .I2(n26513), .O(n26514) );
  MUX2 U28368 ( .A(n26514), .B(img[949]), .S(n28620), .O(n12583) );
  AOI22S U28369 ( .A1(n27065), .A2(img[949]), .B1(n28037), .B2(n30956), .O(
        n26515) );
  ND2S U28370 ( .I1(n26534), .I2(n26515), .O(n26516) );
  AOI22S U28371 ( .A1(n26855), .A2(img[205]), .B1(n24374), .B2(n30957), .O(
        n26517) );
  ND2S U28372 ( .I1(n26534), .I2(n26517), .O(n26518) );
  MUX2 U28373 ( .A(img[181]), .B(n26518), .S(n28626), .O(n13351) );
  AOI22S U28374 ( .A1(n13776), .A2(img[181]), .B1(n28862), .B2(n30958), .O(
        n26519) );
  ND2S U28375 ( .I1(n26534), .I2(n26519), .O(n26520) );
  MUX2 U28376 ( .A(img[205]), .B(n26520), .S(n28629), .O(n13329) );
  AOI22S U28377 ( .A1(n13780), .A2(img[461]), .B1(n28162), .B2(n30959), .O(
        n26521) );
  ND2S U28378 ( .I1(n26534), .I2(n26521), .O(n26522) );
  AOI22S U28379 ( .A1(n13772), .A2(img[437]), .B1(n29407), .B2(n30960), .O(
        n26523) );
  ND2S U28380 ( .I1(n13767), .I2(n26523), .O(n26524) );
  MUX2 U28381 ( .A(n26524), .B(img[461]), .S(n28641), .O(n13073) );
  AOI22S U28382 ( .A1(n13778), .A2(img[1525]), .B1(n28862), .B2(n30961), .O(
        n26525) );
  ND2S U28383 ( .I1(n13767), .I2(n26525), .O(n26526) );
  MUX2 U28384 ( .A(n26526), .B(img[1421]), .S(n28645), .O(n12113) );
  AOI22S U28385 ( .A1(n25062), .A2(n30962), .B1(n26091), .B2(img[1421]), .O(
        n26528) );
  ND2S U28386 ( .I1(n13903), .I2(img[1485]), .O(n26527) );
  ND3S U28387 ( .I1(n26534), .I2(n26528), .I3(n26527), .O(n26529) );
  AOI22S U28388 ( .A1(n28347), .A2(img[1485]), .B1(n28182), .B2(n30963), .O(
        n26530) );
  ND2S U28389 ( .I1(n13767), .I2(n26530), .O(n26531) );
  AOI22S U28390 ( .A1(n25062), .A2(n30964), .B1(n28043), .B2(img[1461]), .O(
        n26533) );
  ND2S U28391 ( .I1(n29258), .I2(img[1525]), .O(n26532) );
  ND3S U28392 ( .I1(n26534), .I2(n26533), .I3(n26532), .O(n26535) );
  MUX2 U28393 ( .A(img[1485]), .B(n26535), .S(n28656), .O(n12049) );
  AOI22S U28394 ( .A1(n28221), .A2(img[845]), .B1(n25468), .B2(n30965), .O(
        n26536) );
  ND2S U28395 ( .I1(n13767), .I2(n26536), .O(n26537) );
  AOI22S U28396 ( .A1(n28221), .A2(img[821]), .B1(n25591), .B2(n30966), .O(
        n26538) );
  ND2S U28397 ( .I1(n13767), .I2(n26538), .O(n26539) );
  MUX2 U28398 ( .A(n26539), .B(img[845]), .S(n28663), .O(n12687) );
  AOI22S U28399 ( .A1(n28221), .A2(img[501]), .B1(n25377), .B2(n30967), .O(
        n26540) );
  ND2S U28400 ( .I1(n13767), .I2(n26540), .O(n26541) );
  MUX2 U28401 ( .A(n26541), .B(img[397]), .S(n29318), .O(n13137) );
  AOI22S U28402 ( .A1(n28221), .A2(img[397]), .B1(n25377), .B2(n30968), .O(
        n26542) );
  ND2S U28403 ( .I1(n13767), .I2(n26542), .O(n26543) );
  MUX2 U28404 ( .A(img[501]), .B(n26543), .S(n29321), .O(n13031) );
  AOI22S U28405 ( .A1(n28412), .A2(img[117]), .B1(n25062), .B2(n30969), .O(
        n26544) );
  ND2S U28406 ( .I1(n13767), .I2(n26544), .O(n26545) );
  AOI22S U28407 ( .A1(n28347), .A2(img[13]), .B1(n28592), .B2(n30970), .O(
        n26546) );
  ND2S U28408 ( .I1(n13767), .I2(n26546), .O(n26547) );
  MUX2 U28409 ( .A(img[117]), .B(n26547), .S(n29536), .O(n13417) );
  AOI22S U28410 ( .A1(n26970), .A2(img[629]), .B1(n13781), .B2(n30971), .O(
        n26548) );
  ND2S U28411 ( .I1(n13767), .I2(n26548), .O(n26549) );
  AOI22S U28412 ( .A1(n28412), .A2(img[525]), .B1(n29530), .B2(n30972), .O(
        n26550) );
  ND2S U28413 ( .I1(n13767), .I2(n26550), .O(n26551) );
  MUX2 U28414 ( .A(n26551), .B(img[629]), .S(n29292), .O(n12905) );
  AOI22S U28415 ( .A1(n27065), .A2(img[1013]), .B1(n29457), .B2(n30973), .O(
        n26552) );
  ND2S U28416 ( .I1(n13767), .I2(n26552), .O(n26553) );
  AOI22S U28417 ( .A1(n24415), .A2(img[909]), .B1(n29242), .B2(n30974), .O(
        n26554) );
  ND2S U28418 ( .I1(n13767), .I2(n26554), .O(n26555) );
  MUX2 U28419 ( .A(img[1013]), .B(n26555), .S(n29303), .O(n12519) );
  AOI22S U28420 ( .A1(n28468), .A2(img[245]), .B1(n23941), .B2(n30975), .O(
        n26556) );
  ND2S U28421 ( .I1(n13767), .I2(n26556), .O(n26557) );
  AOI22S U28422 ( .A1(n26101), .A2(img[141]), .B1(n28614), .B2(n30976), .O(
        n26558) );
  ND2S U28423 ( .I1(n13767), .I2(n26558), .O(n26559) );
  MUX2 U28424 ( .A(img[245]), .B(n26559), .S(n29309), .O(n13287) );
  AOI22S U28425 ( .A1(n13773), .A2(img[373]), .B1(n24374), .B2(n30977), .O(
        n26560) );
  ND2S U28426 ( .I1(n13767), .I2(n26560), .O(n26561) );
  MUX2 U28427 ( .A(n26561), .B(img[269]), .S(n29312), .O(n13263) );
  AOI22S U28428 ( .A1(n25595), .A2(img[269]), .B1(n27511), .B2(n30978), .O(
        n26562) );
  ND2S U28429 ( .I1(n13767), .I2(n26562), .O(n26563) );
  AOI22S U28430 ( .A1(n26101), .A2(img[885]), .B1(n25468), .B2(n30979), .O(
        n26564) );
  ND2S U28431 ( .I1(n13767), .I2(n26564), .O(n26565) );
  INV1S U28432 ( .I(img[885]), .O(n26566) );
  AOI22S U28433 ( .A1(n13777), .A2(img[781]), .B1(n27735), .B2(n26566), .O(
        n26567) );
  ND2S U28434 ( .I1(n13767), .I2(n26567), .O(n26568) );
  MUX2 U28435 ( .A(n26568), .B(img[885]), .S(n29328), .O(n12649) );
  AOI22S U28436 ( .A1(n28221), .A2(img[757]), .B1(n25591), .B2(n30980), .O(
        n26569) );
  ND2S U28437 ( .I1(n13767), .I2(n26569), .O(n26570) );
  AOI22S U28438 ( .A1(n28221), .A2(img[653]), .B1(n29397), .B2(n30981), .O(
        n26571) );
  ND2S U28439 ( .I1(n13767), .I2(n26571), .O(n26572) );
  MUX2 U28440 ( .A(n26572), .B(img[757]), .S(n29334), .O(n12775) );
  AOI22S U28441 ( .A1(n28221), .A2(img[253]), .B1(n24193), .B2(n30982), .O(
        n26573) );
  ND2S U28442 ( .I1(n13767), .I2(n26573), .O(n26574) );
  MUX2 U28443 ( .A(n26574), .B(img[133]), .S(n29402), .O(n13399) );
  AOI22S U28444 ( .A1(n28221), .A2(img[133]), .B1(n13781), .B2(n30983), .O(
        n26575) );
  ND2S U28445 ( .I1(n13767), .I2(n26575), .O(n26576) );
  MUX2 U28446 ( .A(img[253]), .B(n26576), .S(n29405), .O(n13280) );
  AOI22S U28447 ( .A1(n28221), .A2(img[381]), .B1(n29397), .B2(n30984), .O(
        n26577) );
  ND2S U28448 ( .I1(n13767), .I2(n26577), .O(n26578) );
  AOI22S U28449 ( .A1(n28221), .A2(img[261]), .B1(n27511), .B2(n30985), .O(
        n26579) );
  ND2S U28450 ( .I1(n13767), .I2(n26579), .O(n26580) );
  MUX2 U28451 ( .A(img[381]), .B(n26580), .S(n29412), .O(n13151) );
  AOI22S U28452 ( .A1(n29414), .A2(img[637]), .B1(n25591), .B2(n30986), .O(
        n26581) );
  ND2S U28453 ( .I1(n13767), .I2(n26581), .O(n26582) );
  MUX2 U28454 ( .A(n26582), .B(img[517]), .S(n29383), .O(n13017) );
  AOI22S U28455 ( .A1(n29129), .A2(img[517]), .B1(n27511), .B2(n30987), .O(
        n26584) );
  ND2S U28456 ( .I1(n13767), .I2(n26584), .O(n26585) );
  MUX2 U28457 ( .A(n26585), .B(img[637]), .S(n29386), .O(n12895) );
  AOI22S U28458 ( .A1(n13772), .A2(img[125]), .B1(n13781), .B2(n30988), .O(
        n26586) );
  ND2S U28459 ( .I1(n13767), .I2(n26586), .O(n26587) );
  AOI22S U28460 ( .A1(n27957), .A2(img[5]), .B1(n13781), .B2(n30989), .O(
        n26588) );
  ND2S U28461 ( .I1(n13767), .I2(n26588), .O(n26589) );
  MUX2 U28462 ( .A(img[125]), .B(n26589), .S(n29392), .O(n13407) );
  AOI22S U28463 ( .A1(n26101), .A2(img[1021]), .B1(n25062), .B2(n30990), .O(
        n26590) );
  ND2S U28464 ( .I1(n13767), .I2(n26590), .O(n26591) );
  MUX2 U28465 ( .A(img[901]), .B(n26591), .S(n29395), .O(n12631) );
  AOI22S U28466 ( .A1(n28347), .A2(img[901]), .B1(n29457), .B2(n30991), .O(
        n26592) );
  ND2S U28467 ( .I1(n13767), .I2(n26592), .O(n26593) );
  AOI22S U28468 ( .A1(n25595), .A2(img[509]), .B1(n27049), .B2(n30992), .O(
        n26594) );
  ND2S U28469 ( .I1(n13767), .I2(n26594), .O(n26595) );
  INV1S U28470 ( .I(img[509]), .O(n26596) );
  AOI22S U28471 ( .A1(n28347), .A2(img[389]), .B1(n27049), .B2(n26596), .O(
        n26597) );
  ND2S U28472 ( .I1(n13767), .I2(n26597), .O(n26598) );
  MUX2 U28473 ( .A(n26598), .B(img[509]), .S(n29420), .O(n13025) );
  AOI22S U28474 ( .A1(n25595), .A2(img[893]), .B1(n25591), .B2(n30993), .O(
        n26599) );
  ND2S U28475 ( .I1(n13767), .I2(n26599), .O(n26600) );
  INV1S U28476 ( .I(img[893]), .O(n26601) );
  AOI22S U28477 ( .A1(n25810), .A2(img[773]), .B1(n28695), .B2(n26601), .O(
        n26602) );
  ND2S U28478 ( .I1(n13767), .I2(n26602), .O(n26603) );
  MUX2 U28479 ( .A(n26603), .B(img[893]), .S(n29427), .O(n12639) );
  AOI22S U28480 ( .A1(n26101), .A2(img[765]), .B1(n25859), .B2(n30994), .O(
        n26604) );
  ND2S U28481 ( .I1(n13767), .I2(n26604), .O(n26605) );
  AOI22S U28482 ( .A1(n29414), .A2(img[645]), .B1(n13775), .B2(n30995), .O(
        n26606) );
  ND2S U28483 ( .I1(n13767), .I2(n26606), .O(n26607) );
  MUX2 U28484 ( .A(n26607), .B(img[765]), .S(n29433), .O(n12769) );
  AOI22S U28485 ( .A1(n29414), .A2(img[549]), .B1(n25859), .B2(n30996), .O(
        n26608) );
  ND2S U28486 ( .I1(n13767), .I2(n26608), .O(n26609) );
  MUX2 U28487 ( .A(n26609), .B(img[605]), .S(n29478), .O(n12927) );
  AOI22S U28488 ( .A1(n29414), .A2(img[93]), .B1(n24374), .B2(n30997), .O(
        n26610) );
  ND2S U28489 ( .I1(n13767), .I2(n26610), .O(n26611) );
  MUX2 U28490 ( .A(img[37]), .B(n26611), .S(n29342), .O(n13497) );
  AOI22S U28491 ( .A1(n29414), .A2(img[37]), .B1(n27049), .B2(n30998), .O(
        n26612) );
  ND2S U28492 ( .I1(n13767), .I2(n26612), .O(n26613) );
  MUX2 U28493 ( .A(img[93]), .B(n26613), .S(n29339), .O(n13439) );
  AOI22S U28494 ( .A1(n29414), .A2(img[989]), .B1(n25591), .B2(n30999), .O(
        n26614) );
  ND2S U28495 ( .I1(n13767), .I2(n26614), .O(n26615) );
  AOI22S U28496 ( .A1(n27957), .A2(img[933]), .B1(n28343), .B2(n31000), .O(
        n26616) );
  ND2S U28497 ( .I1(n13767), .I2(n26616), .O(n26617) );
  MUX2 U28498 ( .A(img[989]), .B(n26617), .S(n29345), .O(n12545) );
  AOI22S U28499 ( .A1(n27957), .A2(img[221]), .B1(n13775), .B2(n31001), .O(
        n26618) );
  ND2S U28500 ( .I1(n13767), .I2(n26618), .O(n26619) );
  MUX2 U28501 ( .A(img[165]), .B(n26619), .S(n29355), .O(n13367) );
  AOI22S U28502 ( .A1(n27957), .A2(img[165]), .B1(n13775), .B2(n31002), .O(
        n26620) );
  ND2S U28503 ( .I1(n13767), .I2(n26620), .O(n26621) );
  MUX2 U28504 ( .A(img[221]), .B(n26621), .S(n29351), .O(n13313) );
  AOI22S U28505 ( .A1(n27957), .A2(img[349]), .B1(n13775), .B2(n31003), .O(
        n26622) );
  ND2S U28506 ( .I1(n13767), .I2(n26622), .O(n26623) );
  AOI22S U28507 ( .A1(n27957), .A2(img[293]), .B1(n28592), .B2(n31004), .O(
        n26624) );
  ND2S U28508 ( .I1(n13767), .I2(n26624), .O(n26625) );
  MUX2 U28509 ( .A(img[349]), .B(n26625), .S(n29358), .O(n13183) );
  AOI22S U28510 ( .A1(n27957), .A2(img[477]), .B1(n29242), .B2(n31005), .O(
        n26626) );
  ND2S U28511 ( .I1(n13767), .I2(n26626), .O(n26627) );
  MUX2 U28512 ( .A(img[421]), .B(n26627), .S(n29367), .O(n13111) );
  AOI22S U28513 ( .A1(n28347), .A2(img[421]), .B1(n29457), .B2(n31006), .O(
        n26628) );
  ND2S U28514 ( .I1(n13767), .I2(n26628), .O(n26629) );
  MUX2 U28515 ( .A(img[477]), .B(n26629), .S(n29364), .O(n13057) );
  AOI22S U28516 ( .A1(n28347), .A2(img[861]), .B1(n13779), .B2(n31007), .O(
        n26630) );
  ND2S U28517 ( .I1(n13767), .I2(n26630), .O(n26631) );
  MUX2 U28518 ( .A(n26631), .B(img[805]), .S(n29374), .O(n12729) );
  AOI22S U28519 ( .A1(n28347), .A2(img[805]), .B1(n25859), .B2(n31008), .O(
        n26632) );
  ND2S U28520 ( .I1(n13767), .I2(n26632), .O(n26633) );
  AOI22S U28521 ( .A1(n28347), .A2(img[733]), .B1(n24755), .B2(n31009), .O(
        n26634) );
  ND2S U28522 ( .I1(n13767), .I2(n26634), .O(n26635) );
  AOI22S U28523 ( .A1(n29414), .A2(img[677]), .B1(n13781), .B2(n31010), .O(
        n26636) );
  ND2S U28524 ( .I1(n26534), .I2(n26636), .O(n26637) );
  INV1S U28525 ( .I(n29475), .O(n26642) );
  OAI22S U28526 ( .A1(n26639), .A2(n28530), .B1(n13897), .B2(n26638), .O(
        n26640) );
  AOI12HS U28527 ( .B1(n28534), .B2(n29462), .A1(n26640), .O(n26641) );
  OAI12HS U28528 ( .B1(n28536), .B2(n26642), .A1(n26641), .O(n26670) );
  AOI22S U28529 ( .A1(n28552), .A2(A67_shift[137]), .B1(n28553), .B2(
        A67_shift[9]), .O(n26644) );
  ND2S U28530 ( .I1(n28554), .I2(A67_shift[105]), .O(n26643) );
  AOI22S U28531 ( .A1(n28551), .A2(A67_shift[201]), .B1(n28546), .B2(
        A67_shift[169]), .O(n26650) );
  ND2S U28532 ( .I1(A67_shift[233]), .I2(n28547), .O(n26645) );
  ND2S U28533 ( .I1(n28555), .I2(n26645), .O(n26646) );
  AOI12HS U28534 ( .B1(n28550), .B2(A67_shift[73]), .A1(n26646), .O(n26649) );
  INV1S U28535 ( .I(A67_shift[41]), .O(n26647) );
  INV1S U28536 ( .I(A67_shift[185]), .O(n26652) );
  INV1S U28537 ( .I(A67_shift[57]), .O(n26651) );
  OAI22S U28538 ( .A1(n26653), .A2(n26652), .B1(n28544), .B2(n26651), .O(
        n26661) );
  ND2S U28539 ( .I1(n28552), .I2(A67_shift[153]), .O(n26659) );
  AOI22S U28540 ( .A1(n28550), .A2(A67_shift[89]), .B1(n28553), .B2(
        A67_shift[25]), .O(n26658) );
  AOI22S U28541 ( .A1(n28554), .A2(A67_shift[121]), .B1(n28551), .B2(
        A67_shift[217]), .O(n26655) );
  ND2S U28542 ( .I1(A67_shift[249]), .I2(n28547), .O(n26654) );
  ND2S U28543 ( .I1(n26655), .I2(n26654), .O(n26656) );
  NR2 U28544 ( .I1(n26656), .I2(n28555), .O(n26657) );
  OAI22S U28545 ( .A1(n26663), .A2(n26662), .B1(n26661), .B2(n26660), .O(
        n26668) );
  ND2S U28546 ( .I1(n28564), .I2(gray_avg_out[1]), .O(n26666) );
  ND2S U28547 ( .I1(n28565), .I2(gray_weight_out[1]), .O(n26665) );
  ND2S U28548 ( .I1(n28566), .I2(gray_max_out[1]), .O(n26664) );
  AOI22S U28549 ( .A1(n29414), .A2(img[513]), .B1(n13781), .B2(n31011), .O(
        n26671) );
  ND2S U28550 ( .I1(n27156), .I2(n26671), .O(n26672) );
  MUX2 U28551 ( .A(n26672), .B(img[633]), .S(n29386), .O(n12899) );
  AOI22S U28552 ( .A1(n29414), .A2(img[633]), .B1(n29530), .B2(n31012), .O(
        n26673) );
  ND2S U28553 ( .I1(n27156), .I2(n26673), .O(n26674) );
  AOI22S U28554 ( .A1(n29414), .A2(img[1]), .B1(n13779), .B2(n31013), .O(
        n26675) );
  ND2S U28555 ( .I1(n27156), .I2(n26675), .O(n26676) );
  MUX2 U28556 ( .A(img[121]), .B(n26676), .S(n29392), .O(n13411) );
  AOI22S U28557 ( .A1(n29414), .A2(img[121]), .B1(n25591), .B2(n31014), .O(
        n26677) );
  ND2S U28558 ( .I1(n27156), .I2(n26677), .O(n26678) );
  AOI22S U28559 ( .A1(n29414), .A2(img[1217]), .B1(n29530), .B2(n31015), .O(
        n26679) );
  ND2S U28560 ( .I1(n27156), .I2(n26679), .O(n26680) );
  MUX2 U28561 ( .A(img[1209]), .B(n26680), .S(n28821), .O(n12317) );
  BUF12CK U28562 ( .I(n27170), .O(n27156) );
  AOI22S U28563 ( .A1(n28862), .A2(n31016), .B1(n27919), .B2(img[1209]), .O(
        n26682) );
  ND3S U28564 ( .I1(n27156), .I2(n26682), .I3(n26681), .O(n26683) );
  MUX2 U28565 ( .A(img[1217]), .B(n26683), .S(n28818), .O(n12315) );
  AOI22S U28566 ( .A1(n28135), .A2(n31017), .B1(n25444), .B2(img[1153]), .O(
        n26685) );
  ND3S U28567 ( .I1(n27156), .I2(n26685), .I3(n26684), .O(n26686) );
  MUX2 U28568 ( .A(img[1273]), .B(n26686), .S(n28814), .O(n12253) );
  AOI22S U28569 ( .A1(n29414), .A2(img[1273]), .B1(n28614), .B2(n31018), .O(
        n26687) );
  ND2S U28570 ( .I1(n27156), .I2(n26687), .O(n26688) );
  MUX2 U28571 ( .A(img[1153]), .B(n26688), .S(n28810), .O(n12379) );
  AOI22S U28572 ( .A1(n28840), .A2(img[1345]), .B1(n29096), .B2(n31019), .O(
        n26689) );
  ND2S U28573 ( .I1(n27070), .I2(n26689), .O(n26690) );
  AOI22S U28574 ( .A1(n28913), .A2(n31020), .B1(n27919), .B2(img[1337]), .O(
        n26692) );
  ND2S U28575 ( .I1(n13819), .I2(img[1401]), .O(n26691) );
  ND3S U28576 ( .I1(n27156), .I2(n26692), .I3(n26691), .O(n26693) );
  MUX2 U28577 ( .A(img[1345]), .B(n26693), .S(n28832), .O(n12181) );
  AOI22S U28578 ( .A1(n29407), .A2(n31021), .B1(n28254), .B2(img[1281]), .O(
        n26695) );
  ND2S U28579 ( .I1(n13819), .I2(img[1345]), .O(n26694) );
  ND3S U28580 ( .I1(n27156), .I2(n26695), .I3(n26694), .O(n26696) );
  MUX2 U28581 ( .A(img[1401]), .B(n26696), .S(n28828), .O(n12131) );
  AOI22S U28582 ( .A1(n26822), .A2(img[1401]), .B1(n29457), .B2(n31022), .O(
        n26697) );
  ND2S U28583 ( .I1(n27156), .I2(n26697), .O(n26698) );
  AOI22S U28584 ( .A1(n13776), .A2(img[897]), .B1(n29194), .B2(n31023), .O(
        n26699) );
  ND2S U28585 ( .I1(n27070), .I2(n26699), .O(n26700) );
  AOI22S U28586 ( .A1(n29414), .A2(img[1017]), .B1(n25062), .B2(n31024), .O(
        n26701) );
  ND2S U28587 ( .I1(n27156), .I2(n26701), .O(n26702) );
  MUX2 U28588 ( .A(img[897]), .B(n26702), .S(n29395), .O(n12635) );
  AOI22S U28589 ( .A1(n28347), .A2(img[129]), .B1(n24193), .B2(n31025), .O(
        n26703) );
  ND2S U28590 ( .I1(n27156), .I2(n26703), .O(n26704) );
  MUX2 U28591 ( .A(img[249]), .B(n26704), .S(n29405), .O(n13283) );
  AOI22S U28592 ( .A1(n28347), .A2(img[249]), .B1(n28433), .B2(n31026), .O(
        n26705) );
  ND2S U28593 ( .I1(n27156), .I2(n26705), .O(n26706) );
  MUX2 U28594 ( .A(n26706), .B(img[129]), .S(n29402), .O(n13403) );
  AOI22S U28595 ( .A1(n28347), .A2(img[257]), .B1(n29457), .B2(n31027), .O(
        n26707) );
  ND2S U28596 ( .I1(n27070), .I2(n26707), .O(n26708) );
  MUX2 U28597 ( .A(img[377]), .B(n26708), .S(n29412), .O(n13155) );
  AOI22S U28598 ( .A1(n28347), .A2(img[377]), .B1(n25859), .B2(n31028), .O(
        n26709) );
  ND2S U28599 ( .I1(n27070), .I2(n26709), .O(n26710) );
  INV1S U28600 ( .I(img[505]), .O(n26711) );
  AOI22S U28601 ( .A1(n28347), .A2(img[385]), .B1(n28037), .B2(n26711), .O(
        n26712) );
  ND2S U28602 ( .I1(n27156), .I2(n26712), .O(n26713) );
  AOI22S U28603 ( .A1(n28347), .A2(img[505]), .B1(n13781), .B2(n31029), .O(
        n26714) );
  ND2S U28604 ( .I1(n27070), .I2(n26714), .O(n26715) );
  MUX2 U28605 ( .A(n26715), .B(img[385]), .S(n29416), .O(n13147) );
  AOI22S U28606 ( .A1(n28347), .A2(img[1473]), .B1(n25062), .B2(n31030), .O(
        n26716) );
  ND2S U28607 ( .I1(n27070), .I2(n26716), .O(n26717) );
  AOI22S U28608 ( .A1(n28182), .A2(n31031), .B1(n27919), .B2(img[1465]), .O(
        n26719) );
  ND2S U28609 ( .I1(n13819), .I2(img[1529]), .O(n26718) );
  ND3S U28610 ( .I1(n27156), .I2(n26719), .I3(n26718), .O(n26720) );
  MUX2 U28611 ( .A(img[1473]), .B(n26720), .S(n28872), .O(n12059) );
  AOI22S U28612 ( .A1(n25062), .A2(n31032), .B1(n25444), .B2(img[1409]), .O(
        n26722) );
  ND2S U28613 ( .I1(n13819), .I2(img[1473]), .O(n26721) );
  ND3S U28614 ( .I1(n27156), .I2(n26722), .I3(n26721), .O(n26723) );
  AOI22S U28615 ( .A1(n28347), .A2(img[1529]), .B1(n23941), .B2(n31033), .O(
        n26724) );
  ND2S U28616 ( .I1(n27156), .I2(n26724), .O(n26725) );
  MUX2 U28617 ( .A(img[1409]), .B(n26725), .S(n28864), .O(n12123) );
  AOI22S U28618 ( .A1(n28347), .A2(img[769]), .B1(n13781), .B2(n31034), .O(
        n26726) );
  ND2S U28619 ( .I1(n27156), .I2(n26726), .O(n26727) );
  AOI22S U28620 ( .A1(n28347), .A2(img[889]), .B1(n25859), .B2(n31035), .O(
        n26728) );
  ND2S U28621 ( .I1(n27070), .I2(n26728), .O(n26729) );
  MUX2 U28622 ( .A(img[769]), .B(n26729), .S(n29423), .O(n12757) );
  AOI22S U28623 ( .A1(n28347), .A2(img[641]), .B1(n27049), .B2(n31036), .O(
        n26730) );
  ND2S U28624 ( .I1(n27070), .I2(n26730), .O(n26731) );
  AOI22S U28625 ( .A1(n28382), .A2(img[761]), .B1(n28938), .B2(n31037), .O(
        n26732) );
  ND2S U28626 ( .I1(n27156), .I2(n26732), .O(n26733) );
  AOI22S U28627 ( .A1(n27746), .A2(img[1881]), .B1(n25859), .B2(n31038), .O(
        n26734) );
  ND2S U28628 ( .I1(n27156), .I2(n26734), .O(n26735) );
  AOI22S U28629 ( .A1(n29530), .A2(n31039), .B1(n27919), .B2(img[1825]), .O(
        n26737) );
  ND3S U28630 ( .I1(n27070), .I2(n26737), .I3(n26736), .O(n26738) );
  MUX2 U28631 ( .A(img[1881]), .B(n26738), .S(n28896), .O(n11651) );
  AOI22S U28632 ( .A1(n27990), .A2(img[1889]), .B1(n13781), .B2(n31040), .O(
        n26739) );
  ND2S U28633 ( .I1(n27070), .I2(n26739), .O(n26740) );
  MUX2 U28634 ( .A(img[1817]), .B(n26740), .S(n28899), .O(n11715) );
  AOI22S U28635 ( .A1(n29242), .A2(n31041), .B1(n27919), .B2(img[1817]), .O(
        n26742) );
  AOI22S U28636 ( .A1(n13905), .A2(img[1881]), .B1(img[1913]), .B2(n13782), 
        .O(n26741) );
  MUX2 U28637 ( .A(img[1889]), .B(n26743), .S(n28903), .O(n11637) );
  AOI22S U28638 ( .A1(n13773), .A2(img[1857]), .B1(n28182), .B2(n31042), .O(
        n26744) );
  ND2S U28639 ( .I1(n27070), .I2(n26744), .O(n26745) );
  MUX2 U28640 ( .A(img[1849]), .B(n26745), .S(n28919), .O(n11683) );
  AOI22S U28641 ( .A1(n29457), .A2(n31043), .B1(n28254), .B2(img[1849]), .O(
        n26747) );
  ND2S U28642 ( .I1(n13819), .I2(img[1913]), .O(n26746) );
  ND3S U28643 ( .I1(n27156), .I2(n26747), .I3(n26746), .O(n26748) );
  MUX2 U28644 ( .A(img[1857]), .B(n26748), .S(n28916), .O(n11669) );
  AOI22S U28645 ( .A1(n28343), .A2(n31044), .B1(n28254), .B2(img[1793]), .O(
        n26750) );
  AOI22S U28646 ( .A1(n29124), .A2(img[1857]), .B1(img[1889]), .B2(n28908), 
        .O(n26749) );
  ND3S U28647 ( .I1(n27156), .I2(n26750), .I3(n26749), .O(n26751) );
  MUX2 U28648 ( .A(img[1913]), .B(n26751), .S(n28911), .O(n11619) );
  AOI22S U28649 ( .A1(n28083), .A2(img[1913]), .B1(n25859), .B2(n31045), .O(
        n26752) );
  ND2S U28650 ( .I1(n27070), .I2(n26752), .O(n26753) );
  AOI22S U28651 ( .A1(n28083), .A2(img[1753]), .B1(n28862), .B2(n31046), .O(
        n26754) );
  ND2S U28652 ( .I1(n27156), .I2(n26754), .O(n26755) );
  MUX2 U28653 ( .A(n26755), .B(img[1697]), .S(n28922), .O(n11835) );
  AOI22S U28654 ( .A1(n28343), .A2(n31047), .B1(n28254), .B2(img[1697]), .O(
        n26757) );
  ND3S U28655 ( .I1(n27070), .I2(n26757), .I3(n26756), .O(n26758) );
  AOI22S U28656 ( .A1(n27746), .A2(img[1761]), .B1(n13781), .B2(n31048), .O(
        n26759) );
  ND2S U28657 ( .I1(n27156), .I2(n26759), .O(n26760) );
  AOI22S U28658 ( .A1(n28343), .A2(n31049), .B1(n28254), .B2(img[1689]), .O(
        n26762) );
  AOI22S U28659 ( .A1(n29124), .A2(img[1753]), .B1(img[1785]), .B2(n13782), 
        .O(n26761) );
  ND3S U28660 ( .I1(n27070), .I2(n26762), .I3(n26761), .O(n26763) );
  MUX2 U28661 ( .A(img[1761]), .B(n26763), .S(n28933), .O(n11771) );
  AOI22S U28662 ( .A1(n26855), .A2(img[1729]), .B1(n24374), .B2(n31050), .O(
        n26764) );
  ND2S U28663 ( .I1(n27156), .I2(n26764), .O(n26765) );
  MUX2 U28664 ( .A(img[1721]), .B(n26765), .S(n28948), .O(n11805) );
  AOI22S U28665 ( .A1(n25062), .A2(n31051), .B1(n28254), .B2(img[1721]), .O(
        n26767) );
  ND2S U28666 ( .I1(n29124), .I2(img[1785]), .O(n26766) );
  ND3S U28667 ( .I1(n27070), .I2(n26767), .I3(n26766), .O(n26768) );
  MUX2 U28668 ( .A(img[1729]), .B(n26768), .S(n28945), .O(n11803) );
  AOI22S U28669 ( .A1(n25591), .A2(n31052), .B1(n28254), .B2(img[1665]), .O(
        n26770) );
  AOI22S U28670 ( .A1(n29124), .A2(img[1729]), .B1(img[1761]), .B2(n13782), 
        .O(n26769) );
  ND3S U28671 ( .I1(n27070), .I2(n26770), .I3(n26769), .O(n26771) );
  MUX2 U28672 ( .A(img[1785]), .B(n26771), .S(n28941), .O(n11741) );
  AOI22S U28673 ( .A1(n26855), .A2(img[1785]), .B1(n28433), .B2(n31053), .O(
        n26772) );
  ND2S U28674 ( .I1(n27156), .I2(n26772), .O(n26773) );
  AOI22S U28675 ( .A1(n26855), .A2(img[1625]), .B1(n23918), .B2(n31054), .O(
        n26774) );
  ND2S U28676 ( .I1(n27156), .I2(n26774), .O(n26775) );
  MUX2 U28677 ( .A(n26775), .B(img[1569]), .S(n28951), .O(n11957) );
  AOI22S U28678 ( .A1(n28162), .A2(n31055), .B1(n28254), .B2(img[1569]), .O(
        n26777) );
  ND3S U28679 ( .I1(n27070), .I2(n26777), .I3(n26776), .O(n26778) );
  AOI22S U28680 ( .A1(n26855), .A2(img[1633]), .B1(n24755), .B2(n31056), .O(
        n26779) );
  ND2S U28681 ( .I1(n27156), .I2(n26779), .O(n26780) );
  AOI22S U28682 ( .A1(n13779), .A2(n31057), .B1(n28254), .B2(img[1561]), .O(
        n26782) );
  AOI22S U28683 ( .A1(n13770), .A2(img[1625]), .B1(img[1657]), .B2(n13782), 
        .O(n26781) );
  ND3S U28684 ( .I1(n27156), .I2(n26782), .I3(n26781), .O(n26783) );
  MUX2 U28685 ( .A(img[1633]), .B(n26783), .S(n28962), .O(n11899) );
  AOI22S U28686 ( .A1(n28347), .A2(img[1601]), .B1(n28433), .B2(n31058), .O(
        n26784) );
  ND2S U28687 ( .I1(n27070), .I2(n26784), .O(n26785) );
  MUX2 U28688 ( .A(img[1593]), .B(n26785), .S(n28976), .O(n11939) );
  AOI22S U28689 ( .A1(n29096), .A2(n31059), .B1(n28254), .B2(img[1593]), .O(
        n26787) );
  ND3S U28690 ( .I1(n27156), .I2(n26787), .I3(n26786), .O(n26788) );
  MUX2 U28691 ( .A(img[1601]), .B(n26788), .S(n28973), .O(n11925) );
  AOI22S U28692 ( .A1(n29096), .A2(n31060), .B1(n28254), .B2(img[1537]), .O(
        n26790) );
  AOI22S U28693 ( .A1(n13905), .A2(img[1601]), .B1(img[1633]), .B2(n13782), 
        .O(n26789) );
  ND3S U28694 ( .I1(n27070), .I2(n26790), .I3(n26789), .O(n26791) );
  MUX2 U28695 ( .A(img[1657]), .B(n26791), .S(n28969), .O(n11875) );
  AOI22S U28696 ( .A1(n28347), .A2(img[1657]), .B1(n28695), .B2(n31061), .O(
        n26792) );
  ND2S U28697 ( .I1(n27070), .I2(n26792), .O(n26793) );
  AOI22S U28698 ( .A1(n28347), .A2(img[1089]), .B1(n25859), .B2(n31062), .O(
        n26794) );
  ND2S U28699 ( .I1(n27156), .I2(n26794), .O(n26795) );
  AOI22S U28700 ( .A1(n23941), .A2(n31063), .B1(n28254), .B2(img[1081]), .O(
        n26797) );
  ND2S U28701 ( .I1(n13905), .I2(img[1145]), .O(n26796) );
  ND3S U28702 ( .I1(n27156), .I2(n26797), .I3(n26796), .O(n26798) );
  MUX2 U28703 ( .A(img[1089]), .B(n26798), .S(n28987), .O(n12443) );
  AOI22S U28704 ( .A1(n29242), .A2(n31064), .B1(n28069), .B2(img[1025]), .O(
        n26800) );
  ND3S U28705 ( .I1(n27070), .I2(n26800), .I3(n26799), .O(n26801) );
  MUX2 U28706 ( .A(img[1145]), .B(n26801), .S(n28983), .O(n12387) );
  AOI22S U28707 ( .A1(n28347), .A2(img[1145]), .B1(n25062), .B2(n31065), .O(
        n26802) );
  ND2S U28708 ( .I1(n27156), .I2(n26802), .O(n26803) );
  MUX2 U28709 ( .A(img[1025]), .B(n26803), .S(n28979), .O(n12501) );
  AOI22S U28710 ( .A1(n28347), .A2(img[2009]), .B1(n28433), .B2(n31066), .O(
        n26804) );
  ND2S U28711 ( .I1(n27156), .I2(n26804), .O(n26805) );
  MUX2 U28712 ( .A(n26805), .B(img[1953]), .S(n28993), .O(n11579) );
  AOI22S U28713 ( .A1(n28862), .A2(n31067), .B1(n27919), .B2(img[1953]), .O(
        n26807) );
  ND2S U28714 ( .I1(n13820), .I2(img[2017]), .O(n26806) );
  ND3S U28715 ( .I1(n27156), .I2(n26807), .I3(n26806), .O(n26808) );
  AOI22S U28716 ( .A1(n28347), .A2(img[2017]), .B1(n25859), .B2(n31068), .O(
        n26809) );
  ND2S U28717 ( .I1(n27156), .I2(n26809), .O(n26810) );
  MUX2 U28718 ( .A(img[1945]), .B(n26810), .S(n29000), .O(n11581) );
  AOI22S U28719 ( .A1(n28162), .A2(n31069), .B1(n25444), .B2(img[1945]), .O(
        n26812) );
  AOI22S U28720 ( .A1(n13903), .A2(img[2009]), .B1(img[2041]), .B2(n13782), 
        .O(n26811) );
  ND3S U28721 ( .I1(n27156), .I2(n26812), .I3(n26811), .O(n26813) );
  MUX2 U28722 ( .A(img[2017]), .B(n26813), .S(n29004), .O(n11515) );
  AOI22S U28723 ( .A1(n28347), .A2(img[1985]), .B1(n28182), .B2(n31070), .O(
        n26814) );
  ND2S U28724 ( .I1(n27070), .I2(n26814), .O(n26815) );
  MUX2 U28725 ( .A(img[1977]), .B(n26815), .S(n29018), .O(n11549) );
  AOI22S U28726 ( .A1(n13779), .A2(n31071), .B1(n24946), .B2(img[1977]), .O(
        n26817) );
  ND2S U28727 ( .I1(n29124), .I2(img[2041]), .O(n26816) );
  ND3S U28728 ( .I1(n27156), .I2(n26817), .I3(n26816), .O(n26818) );
  MUX2 U28729 ( .A(img[1985]), .B(n26818), .S(n29015), .O(n11547) );
  AOI22S U28730 ( .A1(n28037), .A2(n31072), .B1(n24313), .B2(img[1921]), .O(
        n26820) );
  AOI22S U28731 ( .A1(n13903), .A2(img[1985]), .B1(img[2017]), .B2(n13782), 
        .O(n26819) );
  ND3S U28732 ( .I1(n27156), .I2(n26820), .I3(n26819), .O(n26821) );
  AOI22S U28733 ( .A1(n13780), .A2(img[2041]), .B1(n13779), .B2(n31073), .O(
        n26823) );
  ND2S U28734 ( .I1(n27156), .I2(n26823), .O(n26824) );
  MUX2 U28735 ( .A(img[1921]), .B(n26824), .S(n29007), .O(n11611) );
  AOI22S U28736 ( .A1(n13780), .A2(img[601]), .B1(n13781), .B2(n31074), .O(
        n26825) );
  ND2S U28737 ( .I1(n27156), .I2(n26825), .O(n26826) );
  AOI22S U28738 ( .A1(n13780), .A2(img[33]), .B1(n25468), .B2(n31075), .O(
        n26827) );
  ND2S U28739 ( .I1(n27156), .I2(n26827), .O(n26828) );
  MUX2 U28740 ( .A(img[89]), .B(n26828), .S(n29339), .O(n13443) );
  AOI22S U28741 ( .A1(n13780), .A2(img[89]), .B1(n28592), .B2(n31076), .O(
        n26829) );
  ND2S U28742 ( .I1(n27070), .I2(n26829), .O(n26830) );
  AOI22S U28743 ( .A1(n26855), .A2(img[1249]), .B1(n28075), .B2(n31077), .O(
        n26831) );
  ND2S U28744 ( .I1(n27156), .I2(n26831), .O(n26832) );
  AOI22S U28745 ( .A1(n28075), .A2(n31078), .B1(n24313), .B2(img[1177]), .O(
        n26834) );
  ND2S U28746 ( .I1(n13819), .I2(img[1241]), .O(n26833) );
  ND3S U28747 ( .I1(n27156), .I2(n26834), .I3(n26833), .O(n26835) );
  MUX2 U28748 ( .A(img[1249]), .B(n26835), .S(n29218), .O(n12283) );
  AOI22S U28749 ( .A1(n25062), .A2(n31079), .B1(n24313), .B2(img[1185]), .O(
        n26837) );
  ND2S U28750 ( .I1(n13820), .I2(img[1249]), .O(n26836) );
  ND3S U28751 ( .I1(n27156), .I2(n26837), .I3(n26836), .O(n26838) );
  MUX2 U28752 ( .A(img[1241]), .B(n26838), .S(n29211), .O(n12285) );
  AOI22S U28753 ( .A1(n26855), .A2(img[1241]), .B1(n13775), .B2(n31080), .O(
        n26839) );
  ND2S U28754 ( .I1(n27156), .I2(n26839), .O(n26840) );
  MUX2 U28755 ( .A(n26840), .B(img[1185]), .S(n29207), .O(n12347) );
  AOI22S U28756 ( .A1(n26855), .A2(img[1377]), .B1(n28182), .B2(n31081), .O(
        n26841) );
  ND2S U28757 ( .I1(n27156), .I2(n26841), .O(n26842) );
  MUX2 U28758 ( .A(img[1305]), .B(n26842), .S(n29240), .O(n12227) );
  AOI22S U28759 ( .A1(n29194), .A2(n31082), .B1(n27919), .B2(img[1305]), .O(
        n26844) );
  ND2S U28760 ( .I1(n13904), .I2(img[1369]), .O(n26843) );
  ND3S U28761 ( .I1(n27156), .I2(n26844), .I3(n26843), .O(n26845) );
  MUX2 U28762 ( .A(img[1377]), .B(n26845), .S(n29245), .O(n12149) );
  AOI22S U28763 ( .A1(n28614), .A2(n31083), .B1(n25444), .B2(img[1313]), .O(
        n26847) );
  ND2S U28764 ( .I1(n13905), .I2(img[1377]), .O(n26846) );
  ND3S U28765 ( .I1(n27156), .I2(n26847), .I3(n26846), .O(n26848) );
  MUX2 U28766 ( .A(img[1369]), .B(n26848), .S(n29237), .O(n12163) );
  AOI22S U28767 ( .A1(n26855), .A2(img[1369]), .B1(n25591), .B2(n31084), .O(
        n26849) );
  ND2S U28768 ( .I1(n27156), .I2(n26849), .O(n26850) );
  MUX2 U28769 ( .A(n26850), .B(img[1313]), .S(n29233), .O(n12213) );
  AOI22S U28770 ( .A1(n26855), .A2(img[929]), .B1(n24193), .B2(n31085), .O(
        n26851) );
  ND2S U28771 ( .I1(n27070), .I2(n26851), .O(n26852) );
  MUX2 U28772 ( .A(img[985]), .B(n26852), .S(n29345), .O(n12541) );
  AOI22S U28773 ( .A1(n26855), .A2(img[985]), .B1(n28938), .B2(n31086), .O(
        n26853) );
  ND2S U28774 ( .I1(n27156), .I2(n26853), .O(n26854) );
  AOI22S U28775 ( .A1(n26855), .A2(img[161]), .B1(n28592), .B2(n31087), .O(
        n26856) );
  ND2S U28776 ( .I1(n27156), .I2(n26856), .O(n26857) );
  MUX2 U28777 ( .A(img[217]), .B(n26857), .S(n29351), .O(n13309) );
  AOI22S U28778 ( .A1(n27990), .A2(img[217]), .B1(n25062), .B2(n31088), .O(
        n26858) );
  ND2S U28779 ( .I1(n27156), .I2(n26858), .O(n26859) );
  MUX2 U28780 ( .A(img[161]), .B(n26859), .S(n29355), .O(n13371) );
  AOI22S U28781 ( .A1(n28083), .A2(img[289]), .B1(n25377), .B2(n31089), .O(
        n26860) );
  ND2S U28782 ( .I1(n27156), .I2(n26860), .O(n26861) );
  MUX2 U28783 ( .A(img[345]), .B(n26861), .S(n29358), .O(n13187) );
  AOI22S U28784 ( .A1(n28442), .A2(img[345]), .B1(n13781), .B2(n31090), .O(
        n26862) );
  ND2S U28785 ( .I1(n27070), .I2(n26862), .O(n26863) );
  AOI22S U28786 ( .A1(n28442), .A2(img[417]), .B1(n13775), .B2(n31091), .O(
        n26864) );
  ND2S U28787 ( .I1(n27156), .I2(n26864), .O(n26865) );
  MUX2 U28788 ( .A(img[473]), .B(n26865), .S(n29364), .O(n13053) );
  AOI22S U28789 ( .A1(n13780), .A2(img[473]), .B1(n25468), .B2(n31092), .O(
        n26866) );
  ND2S U28790 ( .I1(n27070), .I2(n26866), .O(n26867) );
  MUX2 U28791 ( .A(img[417]), .B(n26867), .S(n29367), .O(n13115) );
  AOI22S U28792 ( .A1(n13780), .A2(img[1505]), .B1(n29457), .B2(n31093), .O(
        n26868) );
  ND2S U28793 ( .I1(n27070), .I2(n26868), .O(n26869) );
  MUX2 U28794 ( .A(n26869), .B(img[1433]), .S(n29255), .O(n12093) );
  AOI22S U28795 ( .A1(n29194), .A2(n31094), .B1(n28069), .B2(img[1433]), .O(
        n26871) );
  ND3S U28796 ( .I1(n27156), .I2(n26871), .I3(n26870), .O(n26872) );
  MUX2 U28797 ( .A(img[1505]), .B(n26872), .S(n29261), .O(n12027) );
  AOI22S U28798 ( .A1(n28862), .A2(n31095), .B1(n24313), .B2(img[1441]), .O(
        n26874) );
  ND2S U28799 ( .I1(n13820), .I2(img[1505]), .O(n26873) );
  ND3S U28800 ( .I1(n27156), .I2(n26874), .I3(n26873), .O(n26875) );
  AOI22S U28801 ( .A1(n13780), .A2(img[1497]), .B1(n25591), .B2(n31096), .O(
        n26876) );
  ND2S U28802 ( .I1(n27070), .I2(n26876), .O(n26877) );
  MUX2 U28803 ( .A(n26877), .B(img[1441]), .S(n29248), .O(n12091) );
  INV1S U28804 ( .I(img[857]), .O(n26878) );
  AOI22S U28805 ( .A1(n13780), .A2(img[801]), .B1(n28433), .B2(n26878), .O(
        n26879) );
  ND2S U28806 ( .I1(n27156), .I2(n26879), .O(n26880) );
  AOI22S U28807 ( .A1(n13780), .A2(img[857]), .B1(n13781), .B2(n31097), .O(
        n26881) );
  ND2S U28808 ( .I1(n27156), .I2(n26881), .O(n26882) );
  MUX2 U28809 ( .A(n26882), .B(img[801]), .S(n29374), .O(n12725) );
  AOI22S U28810 ( .A1(n13780), .A2(img[673]), .B1(n28695), .B2(n31098), .O(
        n26883) );
  ND2S U28811 ( .I1(n27070), .I2(n26883), .O(n26884) );
  AOI22S U28812 ( .A1(n13780), .A2(img[729]), .B1(n13781), .B2(n31099), .O(
        n26885) );
  ND2S U28813 ( .I1(n27070), .I2(n26885), .O(n26886) );
  AOI22S U28814 ( .A1(n13773), .A2(img[1121]), .B1(n29242), .B2(n31100), .O(
        n26887) );
  ND2S U28815 ( .I1(n27070), .I2(n26887), .O(n26888) );
  AOI22S U28816 ( .A1(n28037), .A2(n31101), .B1(n24313), .B2(img[1049]), .O(
        n26890) );
  ND3S U28817 ( .I1(n27156), .I2(n26890), .I3(n26889), .O(n26891) );
  MUX2 U28818 ( .A(img[1121]), .B(n26891), .S(n29198), .O(n12405) );
  AOI22S U28819 ( .A1(n29194), .A2(n31102), .B1(n24313), .B2(img[1057]), .O(
        n26893) );
  ND3S U28820 ( .I1(n27156), .I2(n26893), .I3(n26892), .O(n26894) );
  MUX2 U28821 ( .A(img[1113]), .B(n26894), .S(n29189), .O(n12419) );
  AOI22S U28822 ( .A1(n27990), .A2(img[1113]), .B1(n28938), .B2(n31103), .O(
        n26895) );
  ND2S U28823 ( .I1(n27070), .I2(n26895), .O(n26896) );
  MUX2 U28824 ( .A(n26896), .B(img[1057]), .S(n29185), .O(n12469) );
  AOI22S U28825 ( .A1(n27746), .A2(img[537]), .B1(n29096), .B2(n31104), .O(
        n26897) );
  ND2S U28826 ( .I1(n27156), .I2(n26897), .O(n26898) );
  MUX2 U28827 ( .A(n26898), .B(img[609]), .S(n29286), .O(n12917) );
  AOI22S U28828 ( .A1(n29414), .A2(img[609]), .B1(n28343), .B2(n31105), .O(
        n26899) );
  ND2S U28829 ( .I1(n27070), .I2(n26899), .O(n26900) );
  AOI22S U28830 ( .A1(n26970), .A2(img[25]), .B1(n25859), .B2(n31106), .O(
        n26901) );
  ND2S U28831 ( .I1(n27070), .I2(n26901), .O(n26902) );
  MUX2 U28832 ( .A(img[97]), .B(n26902), .S(n29280), .O(n13429) );
  AOI22S U28833 ( .A1(n26855), .A2(img[97]), .B1(n28614), .B2(n31107), .O(
        n26903) );
  ND2S U28834 ( .I1(n27070), .I2(n26903), .O(n26904) );
  AOI22S U28835 ( .A1(n28442), .A2(img[921]), .B1(n28037), .B2(n31108), .O(
        n26905) );
  ND2S U28836 ( .I1(n27070), .I2(n26905), .O(n26906) );
  MUX2 U28837 ( .A(img[993]), .B(n26906), .S(n29224), .O(n12539) );
  AOI22S U28838 ( .A1(n27065), .A2(img[993]), .B1(n28182), .B2(n31109), .O(
        n26907) );
  ND2S U28839 ( .I1(n27070), .I2(n26907), .O(n26908) );
  AOI22S U28840 ( .A1(n26970), .A2(img[153]), .B1(n29096), .B2(n31110), .O(
        n26909) );
  ND2S U28841 ( .I1(n27070), .I2(n26909), .O(n26910) );
  MUX2 U28842 ( .A(img[225]), .B(n26910), .S(n29267), .O(n13307) );
  AOI22S U28843 ( .A1(n24415), .A2(img[225]), .B1(n29242), .B2(n31111), .O(
        n26911) );
  ND2S U28844 ( .I1(n27070), .I2(n26911), .O(n26912) );
  MUX2 U28845 ( .A(img[153]), .B(n26912), .S(n29264), .O(n13373) );
  AOI22S U28846 ( .A1(n24415), .A2(img[281]), .B1(n29096), .B2(n31112), .O(
        n26913) );
  ND2S U28847 ( .I1(n27070), .I2(n26913), .O(n26914) );
  MUX2 U28848 ( .A(img[353]), .B(n26914), .S(n29182), .O(n13173) );
  AOI22S U28849 ( .A1(n26970), .A2(img[353]), .B1(n29096), .B2(n31113), .O(
        n26915) );
  ND2S U28850 ( .I1(n27070), .I2(n26915), .O(n26916) );
  AOI22S U28851 ( .A1(n26970), .A2(img[409]), .B1(n25591), .B2(n31114), .O(
        n26917) );
  ND2S U28852 ( .I1(n27070), .I2(n26917), .O(n26918) );
  MUX2 U28853 ( .A(img[481]), .B(n26918), .S(n29273), .O(n13051) );
  AOI22S U28854 ( .A1(n26970), .A2(img[481]), .B1(n13781), .B2(n31115), .O(
        n26919) );
  ND2S U28855 ( .I1(n27070), .I2(n26919), .O(n26920) );
  INV1S U28856 ( .I(img[865]), .O(n26921) );
  AOI22S U28857 ( .A1(n26970), .A2(img[793]), .B1(n13781), .B2(n26921), .O(
        n26922) );
  ND2S U28858 ( .I1(n27156), .I2(n26922), .O(n26923) );
  AOI22S U28859 ( .A1(n28083), .A2(img[865]), .B1(n13781), .B2(n31116), .O(
        n26924) );
  ND2S U28860 ( .I1(n27070), .I2(n26924), .O(n26925) );
  MUX2 U28861 ( .A(img[793]), .B(n26925), .S(n29227), .O(n12739) );
  AOI22S U28862 ( .A1(n28382), .A2(img[665]), .B1(n13781), .B2(n31117), .O(
        n26926) );
  ND2S U28863 ( .I1(n27070), .I2(n26926), .O(n26927) );
  AOI22S U28864 ( .A1(n26822), .A2(img[737]), .B1(n13781), .B2(n31118), .O(
        n26928) );
  ND2S U28865 ( .I1(n27070), .I2(n26928), .O(n26929) );
  AOI22S U28866 ( .A1(n26822), .A2(img[593]), .B1(n13781), .B2(n31119), .O(
        n26930) );
  ND2S U28867 ( .I1(n27070), .I2(n26930), .O(n26931) );
  MUX2 U28868 ( .A(n26931), .B(img[553]), .S(n29439), .O(n12979) );
  AOI22S U28869 ( .A1(n28382), .A2(img[553]), .B1(n13781), .B2(n31120), .O(
        n26932) );
  ND2S U28870 ( .I1(n27156), .I2(n26932), .O(n26933) );
  MUX2 U28871 ( .A(n26933), .B(img[593]), .S(n29133), .O(n12933) );
  AOI22S U28872 ( .A1(n29414), .A2(img[81]), .B1(n13781), .B2(n31121), .O(
        n26934) );
  ND2S U28873 ( .I1(n27070), .I2(n26934), .O(n26935) );
  MUX2 U28874 ( .A(img[41]), .B(n26935), .S(n29136), .O(n13491) );
  AOI22S U28875 ( .A1(n27746), .A2(img[41]), .B1(n13781), .B2(n31122), .O(
        n26936) );
  ND2S U28876 ( .I1(n27070), .I2(n26936), .O(n26937) );
  AOI22S U28877 ( .A1(n29435), .A2(img[1257]), .B1(n25062), .B2(n31123), .O(
        n26938) );
  ND2S U28878 ( .I1(n27070), .I2(n26938), .O(n26939) );
  MUX2 U28879 ( .A(img[1169]), .B(n26939), .S(n29040), .O(n12363) );
  AOI22S U28880 ( .A1(n27735), .A2(n31124), .B1(n24313), .B2(img[1169]), .O(
        n26941) );
  ND3S U28881 ( .I1(n27070), .I2(n26941), .I3(n26940), .O(n26942) );
  MUX2 U28882 ( .A(img[1257]), .B(n26942), .S(n29044), .O(n12269) );
  AOI22S U28883 ( .A1(n28347), .A2(img[1233]), .B1(n28862), .B2(n31125), .O(
        n26943) );
  ND2S U28884 ( .I1(n27070), .I2(n26943), .O(n26944) );
  AOI22S U28885 ( .A1(n24193), .A2(n31126), .B1(n24313), .B2(img[1193]), .O(
        n26946) );
  ND2S U28886 ( .I1(n13819), .I2(img[1257]), .O(n26945) );
  ND3S U28887 ( .I1(n27156), .I2(n26946), .I3(n26945), .O(n26947) );
  MUX2 U28888 ( .A(img[1233]), .B(n26947), .S(n29037), .O(n12299) );
  AOI22S U28889 ( .A1(n26970), .A2(img[1385]), .B1(n28135), .B2(n31127), .O(
        n26948) );
  ND2S U28890 ( .I1(n27070), .I2(n26948), .O(n26949) );
  MUX2 U28891 ( .A(n26949), .B(img[1297]), .S(n29054), .O(n12229) );
  AOI22S U28892 ( .A1(n25377), .A2(n31128), .B1(n24313), .B2(img[1297]), .O(
        n26951) );
  ND3S U28893 ( .I1(n27070), .I2(n26951), .I3(n26950), .O(n26952) );
  MUX2 U28894 ( .A(img[1385]), .B(n26952), .S(n29058), .O(n12147) );
  AOI22S U28895 ( .A1(n28442), .A2(img[1361]), .B1(n28614), .B2(n31129), .O(
        n26953) );
  ND2S U28896 ( .I1(n27156), .I2(n26953), .O(n26954) );
  AOI22S U28897 ( .A1(n29096), .A2(n31130), .B1(n24313), .B2(img[1321]), .O(
        n26956) );
  ND3S U28898 ( .I1(n27156), .I2(n26956), .I3(n26955), .O(n26957) );
  MUX2 U28899 ( .A(img[1361]), .B(n26957), .S(n29051), .O(n12165) );
  AOI22S U28900 ( .A1(n26970), .A2(img[977]), .B1(n28182), .B2(n31131), .O(
        n26958) );
  ND2S U28901 ( .I1(n27156), .I2(n26958), .O(n26959) );
  MUX2 U28902 ( .A(n26959), .B(img[937]), .S(n29142), .O(n12591) );
  AOI22S U28903 ( .A1(n26970), .A2(img[937]), .B1(n28182), .B2(n31132), .O(
        n26960) );
  ND2S U28904 ( .I1(n27156), .I2(n26960), .O(n26961) );
  AOI22S U28905 ( .A1(n26970), .A2(img[209]), .B1(n29242), .B2(n31133), .O(
        n26962) );
  ND2S U28906 ( .I1(n27156), .I2(n26962), .O(n26963) );
  MUX2 U28907 ( .A(img[169]), .B(n26963), .S(n29148), .O(n13357) );
  AOI22S U28908 ( .A1(n26970), .A2(img[169]), .B1(n28182), .B2(n31134), .O(
        n26964) );
  ND2S U28909 ( .I1(n27070), .I2(n26964), .O(n26965) );
  MUX2 U28910 ( .A(img[209]), .B(n26965), .S(n29151), .O(n13323) );
  AOI22S U28911 ( .A1(n26970), .A2(img[337]), .B1(n24755), .B2(n31135), .O(
        n26966) );
  ND2S U28912 ( .I1(n27156), .I2(n26966), .O(n26967) );
  AOI22S U28913 ( .A1(n26970), .A2(img[297]), .B1(n28162), .B2(n31136), .O(
        n26968) );
  ND2S U28914 ( .I1(n27156), .I2(n26968), .O(n26969) );
  MUX2 U28915 ( .A(img[337]), .B(n26969), .S(n29157), .O(n13189) );
  AOI22S U28916 ( .A1(n26970), .A2(img[465]), .B1(n28162), .B2(n31137), .O(
        n26971) );
  ND2S U28917 ( .I1(n27156), .I2(n26971), .O(n26972) );
  AOI22S U28918 ( .A1(n27065), .A2(img[425]), .B1(n28913), .B2(n31138), .O(
        n26973) );
  ND2S U28919 ( .I1(n27070), .I2(n26973), .O(n26974) );
  MUX2 U28920 ( .A(img[465]), .B(n26974), .S(n29163), .O(n13067) );
  AOI22S U28921 ( .A1(n27065), .A2(img[1513]), .B1(n29457), .B2(n31139), .O(
        n26975) );
  ND2S U28922 ( .I1(n27156), .I2(n26975), .O(n26976) );
  AOI22S U28923 ( .A1(n29242), .A2(n31140), .B1(n24313), .B2(img[1425]), .O(
        n26978) );
  ND3S U28924 ( .I1(n27156), .I2(n26978), .I3(n26977), .O(n26979) );
  MUX2 U28925 ( .A(img[1513]), .B(n26979), .S(n29099), .O(n12013) );
  AOI22S U28926 ( .A1(n27065), .A2(img[1489]), .B1(n28913), .B2(n31141), .O(
        n26980) );
  ND2S U28927 ( .I1(n27156), .I2(n26980), .O(n26981) );
  MUX2 U28928 ( .A(n26981), .B(img[1449]), .S(n29087), .O(n12077) );
  AOI22S U28929 ( .A1(n28135), .A2(n31142), .B1(n24313), .B2(img[1449]), .O(
        n26983) );
  ND2S U28930 ( .I1(n13819), .I2(img[1513]), .O(n26982) );
  AOI22S U28931 ( .A1(n27065), .A2(img[849]), .B1(n29407), .B2(n31143), .O(
        n26985) );
  ND2S U28932 ( .I1(n27070), .I2(n26985), .O(n26986) );
  MUX2 U28933 ( .A(n26986), .B(img[809]), .S(n29166), .O(n12723) );
  INV1S U28934 ( .I(img[849]), .O(n26987) );
  AOI22S U28935 ( .A1(n27065), .A2(img[809]), .B1(n29194), .B2(n26987), .O(
        n26988) );
  ND2S U28936 ( .I1(n27070), .I2(n26988), .O(n26989) );
  AOI22S U28937 ( .A1(n24415), .A2(img[721]), .B1(n24755), .B2(n31144), .O(
        n26990) );
  ND2S U28938 ( .I1(n27070), .I2(n26990), .O(n26991) );
  AOI22S U28939 ( .A1(n28347), .A2(img[681]), .B1(n28182), .B2(n31145), .O(
        n26992) );
  ND2S U28940 ( .I1(n27156), .I2(n26992), .O(n26993) );
  AOI22S U28941 ( .A1(n28347), .A2(img[1865]), .B1(n28162), .B2(n31146), .O(
        n26994) );
  ND2S U28942 ( .I1(n27070), .I2(n26994), .O(n26995) );
  MUX2 U28943 ( .A(n26995), .B(img[1841]), .S(n28693), .O(n11685) );
  AOI22S U28944 ( .A1(n25591), .A2(n31147), .B1(n24313), .B2(img[1841]), .O(
        n26997) );
  ND3S U28945 ( .I1(n27156), .I2(n26997), .I3(n26996), .O(n26998) );
  MUX2 U28946 ( .A(img[1865]), .B(n26998), .S(n28698), .O(n11667) );
  AOI22S U28947 ( .A1(n28106), .A2(img[1905]), .B1(n25859), .B2(n31148), .O(
        n26999) );
  ND2S U28948 ( .I1(n27156), .I2(n26999), .O(n27000) );
  AOI22S U28949 ( .A1(n29096), .A2(n31149), .B1(n24313), .B2(img[1801]), .O(
        n27002) );
  AOI22S U28950 ( .A1(n13903), .A2(img[1865]), .B1(img[1897]), .B2(n13782), 
        .O(n27001) );
  ND3S U28951 ( .I1(n27156), .I2(n27002), .I3(n27001), .O(n27003) );
  MUX2 U28952 ( .A(img[1905]), .B(n27003), .S(n28690), .O(n11621) );
  AOI22S U28953 ( .A1(n26855), .A2(img[1897]), .B1(n13781), .B2(n31150), .O(
        n27004) );
  ND2S U28954 ( .I1(n27156), .I2(n27004), .O(n27005) );
  MUX2 U28955 ( .A(n27005), .B(img[1809]), .S(n28679), .O(n11717) );
  AOI22S U28956 ( .A1(n28913), .A2(n31151), .B1(n24313), .B2(img[1809]), .O(
        n27007) );
  AOI22S U28957 ( .A1(n29258), .A2(img[1873]), .B1(img[1905]), .B2(n13782), 
        .O(n27006) );
  ND3S U28958 ( .I1(n27156), .I2(n27007), .I3(n27006), .O(n27008) );
  MUX2 U28959 ( .A(img[1897]), .B(n27008), .S(n28683), .O(n11635) );
  AOI22S U28960 ( .A1(n24415), .A2(img[1873]), .B1(n28938), .B2(n31152), .O(
        n27009) );
  ND2S U28961 ( .I1(n27156), .I2(n27009), .O(n27010) );
  MUX2 U28962 ( .A(n27010), .B(img[1833]), .S(n28672), .O(n11699) );
  AOI22S U28963 ( .A1(n29242), .A2(n31153), .B1(n28069), .B2(img[1833]), .O(
        n27012) );
  ND2S U28964 ( .I1(n13819), .I2(img[1897]), .O(n27011) );
  ND3S U28965 ( .I1(n27156), .I2(n27012), .I3(n27011), .O(n27013) );
  MUX2 U28966 ( .A(img[1873]), .B(n27013), .S(n28676), .O(n11653) );
  AOI22S U28967 ( .A1(n28347), .A2(img[1737]), .B1(n25859), .B2(n31154), .O(
        n27014) );
  ND2S U28968 ( .I1(n27070), .I2(n27014), .O(n27015) );
  MUX2 U28969 ( .A(n27015), .B(img[1713]), .S(n28722), .O(n11819) );
  AOI22S U28970 ( .A1(n28862), .A2(n31155), .B1(n26504), .B2(img[1713]), .O(
        n27017) );
  ND3S U28971 ( .I1(n27156), .I2(n27017), .I3(n27016), .O(n27018) );
  MUX2 U28972 ( .A(img[1737]), .B(n27018), .S(n28726), .O(n11789) );
  AOI22S U28973 ( .A1(n28347), .A2(img[1777]), .B1(n27049), .B2(n31156), .O(
        n27019) );
  ND2S U28974 ( .I1(n27156), .I2(n27019), .O(n27020) );
  AOI22S U28975 ( .A1(n28913), .A2(n31157), .B1(n29257), .B2(img[1673]), .O(
        n27022) );
  AOI22S U28976 ( .A1(n13904), .A2(img[1737]), .B1(img[1769]), .B2(n13782), 
        .O(n27021) );
  ND3S U28977 ( .I1(n27156), .I2(n27022), .I3(n27021), .O(n27023) );
  MUX2 U28978 ( .A(img[1777]), .B(n27023), .S(n28719), .O(n11755) );
  AOI22S U28979 ( .A1(n28347), .A2(img[1769]), .B1(n29242), .B2(n31158), .O(
        n27024) );
  ND2S U28980 ( .I1(n27156), .I2(n27024), .O(n27025) );
  AOI22S U28981 ( .A1(n13781), .A2(n31159), .B1(n26091), .B2(img[1681]), .O(
        n27027) );
  AOI22S U28982 ( .A1(n13903), .A2(img[1745]), .B1(img[1777]), .B2(n13782), 
        .O(n27026) );
  ND3 U28983 ( .I1(n27170), .I2(n27027), .I3(n27026), .O(n27028) );
  AOI22S U28984 ( .A1(n28442), .A2(img[1745]), .B1(n28913), .B2(n31160), .O(
        n27029) );
  ND2S U28985 ( .I1(n27156), .I2(n27029), .O(n27030) );
  AOI22S U28986 ( .A1(n29242), .A2(n31161), .B1(n24946), .B2(img[1705]), .O(
        n27032) );
  ND2S U28987 ( .I1(n13901), .I2(img[1769]), .O(n27031) );
  ND3S U28988 ( .I1(n27156), .I2(n27032), .I3(n27031), .O(n27033) );
  MUX2 U28989 ( .A(img[1745]), .B(n27033), .S(n28705), .O(n11787) );
  AOI22S U28990 ( .A1(n27065), .A2(img[1609]), .B1(n28695), .B2(n31162), .O(
        n27034) );
  ND2S U28991 ( .I1(n27156), .I2(n27034), .O(n27035) );
  AOI22S U28992 ( .A1(n25591), .A2(n31163), .B1(n28069), .B2(img[1585]), .O(
        n27037) );
  ND2S U28993 ( .I1(n29124), .I2(img[1649]), .O(n27036) );
  ND3S U28994 ( .I1(n27156), .I2(n27037), .I3(n27036), .O(n27038) );
  MUX2 U28995 ( .A(img[1609]), .B(n27038), .S(n28754), .O(n11923) );
  AOI22S U28996 ( .A1(n27065), .A2(img[1649]), .B1(n29407), .B2(n31164), .O(
        n27039) );
  ND2S U28997 ( .I1(n27156), .I2(n27039), .O(n27040) );
  AOI22S U28998 ( .A1(n28913), .A2(n31165), .B1(n25444), .B2(img[1545]), .O(
        n27042) );
  AOI22S U28999 ( .A1(n13905), .A2(img[1609]), .B1(img[1641]), .B2(n13782), 
        .O(n27041) );
  ND3S U29000 ( .I1(n27156), .I2(n27042), .I3(n27041), .O(n27043) );
  MUX2 U29001 ( .A(img[1649]), .B(n27043), .S(n28747), .O(n11877) );
  AOI22S U29002 ( .A1(n27065), .A2(img[1641]), .B1(n25591), .B2(n31166), .O(
        n27044) );
  ND2S U29003 ( .I1(n27156), .I2(n27044), .O(n27045) );
  MUX2 U29004 ( .A(n27045), .B(img[1553]), .S(n28736), .O(n11973) );
  AOI22S U29005 ( .A1(n13781), .A2(n31167), .B1(n29257), .B2(img[1553]), .O(
        n27047) );
  AOI22S U29006 ( .A1(n13905), .A2(img[1617]), .B1(img[1649]), .B2(n13782), 
        .O(n27046) );
  ND3S U29007 ( .I1(n27156), .I2(n27047), .I3(n27046), .O(n27048) );
  MUX2 U29008 ( .A(img[1641]), .B(n27048), .S(n28740), .O(n11891) );
  AOI22S U29009 ( .A1(n27065), .A2(img[1617]), .B1(n27049), .B2(n31168), .O(
        n27050) );
  ND2S U29010 ( .I1(n27156), .I2(n27050), .O(n27051) );
  MUX2 U29011 ( .A(n27051), .B(img[1577]), .S(n28729), .O(n11955) );
  AOI22S U29012 ( .A1(n29242), .A2(n31169), .B1(n26504), .B2(img[1577]), .O(
        n27053) );
  ND3S U29013 ( .I1(n27156), .I2(n27053), .I3(n27052), .O(n27054) );
  MUX2 U29014 ( .A(img[1617]), .B(n27054), .S(n28733), .O(n11909) );
  AOI22S U29015 ( .A1(n27065), .A2(img[1129]), .B1(n24193), .B2(n31170), .O(
        n27055) );
  ND2S U29016 ( .I1(n27156), .I2(n27055), .O(n27056) );
  AOI22S U29017 ( .A1(n25377), .A2(n31171), .B1(n24434), .B2(img[1041]), .O(
        n27058) );
  ND2S U29018 ( .I1(n13820), .I2(img[1105]), .O(n27057) );
  ND3S U29019 ( .I1(n27156), .I2(n27058), .I3(n27057), .O(n27059) );
  MUX2 U29020 ( .A(img[1129]), .B(n27059), .S(n29127), .O(n12403) );
  AOI22S U29021 ( .A1(n27065), .A2(img[1105]), .B1(n28135), .B2(n31172), .O(
        n27060) );
  ND2S U29022 ( .I1(n27156), .I2(n27060), .O(n27061) );
  MUX2 U29023 ( .A(n27061), .B(img[1065]), .S(n29115), .O(n12467) );
  AOI22S U29024 ( .A1(n28343), .A2(n31173), .B1(n24946), .B2(img[1065]), .O(
        n27063) );
  ND3S U29025 ( .I1(n27156), .I2(n27063), .I3(n27062), .O(n27064) );
  MUX2 U29026 ( .A(img[1105]), .B(n27064), .S(n29119), .O(n12421) );
  AOI22S U29027 ( .A1(n27065), .A2(img[1993]), .B1(n29194), .B2(n31174), .O(
        n27066) );
  ND2S U29028 ( .I1(n27156), .I2(n27066), .O(n27067) );
  MUX2 U29029 ( .A(n27067), .B(img[1969]), .S(n28792), .O(n11563) );
  AOI22S U29030 ( .A1(n28938), .A2(n31175), .B1(n28069), .B2(img[1969]), .O(
        n27069) );
  ND3S U29031 ( .I1(n27070), .I2(n27069), .I3(n27068), .O(n27071) );
  MUX2 U29032 ( .A(img[1993]), .B(n27071), .S(n28796), .O(n11533) );
  AOI22S U29033 ( .A1(n28106), .A2(img[2033]), .B1(n27443), .B2(n31176), .O(
        n27072) );
  ND2S U29034 ( .I1(n27156), .I2(n27072), .O(n27073) );
  MUX2 U29035 ( .A(img[1929]), .B(n27073), .S(n28785), .O(n11597) );
  AOI22S U29036 ( .A1(n28862), .A2(n31177), .B1(n28069), .B2(img[1929]), .O(
        n27075) );
  AOI22S U29037 ( .A1(n13820), .A2(img[1993]), .B1(img[2025]), .B2(n13782), 
        .O(n27074) );
  ND3S U29038 ( .I1(n27156), .I2(n27075), .I3(n27074), .O(n27076) );
  MUX2 U29039 ( .A(img[2033]), .B(n27076), .S(n28789), .O(n11499) );
  AOI22S U29040 ( .A1(n28347), .A2(img[2025]), .B1(n28862), .B2(n31178), .O(
        n27077) );
  ND2S U29041 ( .I1(n27156), .I2(n27077), .O(n27078) );
  MUX2 U29042 ( .A(n27078), .B(img[1937]), .S(n28778), .O(n11595) );
  AOI22S U29043 ( .A1(n28862), .A2(n31179), .B1(n28069), .B2(img[1937]), .O(
        n27080) );
  AOI22S U29044 ( .A1(n13905), .A2(img[2001]), .B1(img[2033]), .B2(n13782), 
        .O(n27079) );
  ND3S U29045 ( .I1(n27156), .I2(n27080), .I3(n27079), .O(n27081) );
  MUX2 U29046 ( .A(img[2025]), .B(n27081), .S(n28782), .O(n11501) );
  AOI22S U29047 ( .A1(n27065), .A2(img[2001]), .B1(n25591), .B2(n31180), .O(
        n27082) );
  ND2S U29048 ( .I1(n27156), .I2(n27082), .O(n27083) );
  MUX2 U29049 ( .A(n27083), .B(img[1961]), .S(n28771), .O(n11565) );
  AOI22S U29050 ( .A1(n24193), .A2(n31181), .B1(n28069), .B2(img[1961]), .O(
        n27085) );
  ND3S U29051 ( .I1(n27156), .I2(n27085), .I3(n27084), .O(n27086) );
  MUX2 U29052 ( .A(img[2001]), .B(n27086), .S(n28775), .O(n11531) );
  AOI22S U29053 ( .A1(n25595), .A2(img[1225]), .B1(n24193), .B2(n31182), .O(
        n27087) );
  ND2S U29054 ( .I1(n27070), .I2(n27087), .O(n27088) );
  AOI22S U29055 ( .A1(n25062), .A2(n31183), .B1(n28069), .B2(img[1201]), .O(
        n27090) );
  ND2S U29056 ( .I1(n29124), .I2(img[1265]), .O(n27089) );
  ND3S U29057 ( .I1(n27156), .I2(n27090), .I3(n27089), .O(n27091) );
  MUX2 U29058 ( .A(img[1225]), .B(n27091), .S(n28602), .O(n12301) );
  AOI22S U29059 ( .A1(n27990), .A2(img[1265]), .B1(n25377), .B2(n31184), .O(
        n27092) );
  ND2S U29060 ( .I1(n27156), .I2(n27092), .O(n27093) );
  AOI22S U29061 ( .A1(n28075), .A2(n31185), .B1(n28069), .B2(img[1161]), .O(
        n27095) );
  ND2S U29062 ( .I1(n29124), .I2(img[1225]), .O(n27094) );
  ND3S U29063 ( .I1(n27156), .I2(n27095), .I3(n27094), .O(n27096) );
  MUX2 U29064 ( .A(img[1265]), .B(n27096), .S(n28595), .O(n12267) );
  AOI22S U29065 ( .A1(n29414), .A2(img[881]), .B1(n23918), .B2(n31186), .O(
        n27097) );
  ND2S U29066 ( .I1(n27156), .I2(n27097), .O(n27098) );
  MUX2 U29067 ( .A(img[777]), .B(n27098), .S(n29324), .O(n12755) );
  INV1S U29068 ( .I(img[881]), .O(n27099) );
  AOI22S U29069 ( .A1(n27746), .A2(img[777]), .B1(n28695), .B2(n27099), .O(
        n27100) );
  ND2S U29070 ( .I1(n27156), .I2(n27100), .O(n27101) );
  AOI22S U29071 ( .A1(n13777), .A2(img[625]), .B1(n13779), .B2(n31187), .O(
        n27102) );
  ND2S U29072 ( .I1(n27156), .I2(n27102), .O(n27103) );
  AOI22S U29073 ( .A1(n13776), .A2(img[521]), .B1(n23941), .B2(n31188), .O(
        n27104) );
  ND2S U29074 ( .I1(n27156), .I2(n27104), .O(n27105) );
  MUX2 U29075 ( .A(n27105), .B(img[625]), .S(n29292), .O(n12901) );
  AOI22S U29076 ( .A1(n28083), .A2(img[113]), .B1(n29530), .B2(n31189), .O(
        n27106) );
  ND2S U29077 ( .I1(n27156), .I2(n27106), .O(n27107) );
  MUX2 U29078 ( .A(n27107), .B(img[9]), .S(n29295), .O(n13523) );
  AOI22S U29079 ( .A1(n26855), .A2(img[9]), .B1(n25377), .B2(n31190), .O(
        n27108) );
  ND2S U29080 ( .I1(n27156), .I2(n27108), .O(n27109) );
  AOI22S U29081 ( .A1(n24415), .A2(img[1353]), .B1(n23918), .B2(n31191), .O(
        n27111) );
  ND2S U29082 ( .I1(n27156), .I2(n27111), .O(n27112) );
  MUX2 U29083 ( .A(n27112), .B(img[1329]), .S(n28612), .O(n12197) );
  AOI22S U29084 ( .A1(n13779), .A2(n31192), .B1(n28069), .B2(img[1329]), .O(
        n27114) );
  ND2S U29085 ( .I1(n29124), .I2(img[1393]), .O(n27113) );
  ND3S U29086 ( .I1(n27156), .I2(n27114), .I3(n27113), .O(n27115) );
  MUX2 U29087 ( .A(img[1353]), .B(n27115), .S(n28617), .O(n12179) );
  AOI22S U29088 ( .A1(n29435), .A2(img[1393]), .B1(n28695), .B2(n31193), .O(
        n27116) );
  ND2S U29089 ( .I1(n27070), .I2(n27116), .O(n27117) );
  MUX2 U29090 ( .A(img[1289]), .B(n27117), .S(n28605), .O(n12243) );
  AOI22S U29091 ( .A1(n29096), .A2(n31194), .B1(n28069), .B2(img[1289]), .O(
        n27119) );
  ND3S U29092 ( .I1(n27156), .I2(n27119), .I3(n27118), .O(n27120) );
  MUX2 U29093 ( .A(img[1393]), .B(n27120), .S(n28609), .O(n12133) );
  AOI22S U29094 ( .A1(n28442), .A2(img[241]), .B1(n25591), .B2(n31195), .O(
        n27121) );
  ND2S U29095 ( .I1(n27156), .I2(n27121), .O(n27122) );
  AOI22S U29096 ( .A1(n13773), .A2(img[137]), .B1(n28862), .B2(n31196), .O(
        n27123) );
  ND2S U29097 ( .I1(n27156), .I2(n27123), .O(n27124) );
  MUX2 U29098 ( .A(img[241]), .B(n27124), .S(n29309), .O(n13291) );
  AOI22S U29099 ( .A1(n28442), .A2(img[369]), .B1(n28862), .B2(n31197), .O(
        n27125) );
  ND2S U29100 ( .I1(n27156), .I2(n27125), .O(n27126) );
  MUX2 U29101 ( .A(n27126), .B(img[265]), .S(n29312), .O(n13267) );
  AOI22S U29102 ( .A1(n29435), .A2(img[265]), .B1(n27511), .B2(n31198), .O(
        n27127) );
  ND2S U29103 ( .I1(n27070), .I2(n27127), .O(n27128) );
  AOI22S U29104 ( .A1(n29072), .A2(img[497]), .B1(n24755), .B2(n31199), .O(
        n27129) );
  ND2S U29105 ( .I1(n27156), .I2(n27129), .O(n27130) );
  MUX2 U29106 ( .A(n27130), .B(img[393]), .S(n29318), .O(n13133) );
  AOI22S U29107 ( .A1(n28106), .A2(img[393]), .B1(n27511), .B2(n31200), .O(
        n27131) );
  ND2S U29108 ( .I1(n27156), .I2(n27131), .O(n27132) );
  MUX2 U29109 ( .A(img[497]), .B(n27132), .S(n29321), .O(n13035) );
  AOI22S U29110 ( .A1(n24415), .A2(img[1481]), .B1(n27735), .B2(n31201), .O(
        n27133) );
  ND2S U29111 ( .I1(n27156), .I2(n27133), .O(n27134) );
  AOI22S U29112 ( .A1(n28343), .A2(n31202), .B1(n28069), .B2(img[1457]), .O(
        n27136) );
  ND2S U29113 ( .I1(n13820), .I2(img[1521]), .O(n27135) );
  ND3S U29114 ( .I1(n27156), .I2(n27136), .I3(n27135), .O(n27137) );
  MUX2 U29115 ( .A(img[1481]), .B(n27137), .S(n28656), .O(n12045) );
  AOI22S U29116 ( .A1(n26970), .A2(img[1521]), .B1(n27735), .B2(n31203), .O(
        n27138) );
  ND2S U29117 ( .I1(n27070), .I2(n27138), .O(n27139) );
  MUX2 U29118 ( .A(n27139), .B(img[1417]), .S(n28645), .O(n12109) );
  AOI22S U29119 ( .A1(n28037), .A2(n31204), .B1(n28069), .B2(img[1417]), .O(
        n27141) );
  ND3S U29120 ( .I1(n27156), .I2(n27141), .I3(n27140), .O(n27142) );
  AOI22S U29121 ( .A1(n26822), .A2(img[753]), .B1(n23941), .B2(n31205), .O(
        n27143) );
  ND2S U29122 ( .I1(n27070), .I2(n27143), .O(n27144) );
  MUX2 U29123 ( .A(img[649]), .B(n27144), .S(n29331), .O(n12877) );
  AOI22S U29124 ( .A1(n13780), .A2(img[649]), .B1(n25591), .B2(n31206), .O(
        n27145) );
  ND2S U29125 ( .I1(n27156), .I2(n27145), .O(n27146) );
  AOI22S U29126 ( .A1(n13778), .A2(img[1097]), .B1(n13781), .B2(n31207), .O(
        n27147) );
  ND2S U29127 ( .I1(n27070), .I2(n27147), .O(n27148) );
  MUX2 U29128 ( .A(n27148), .B(img[1073]), .S(n28764), .O(n12453) );
  AOI22S U29129 ( .A1(n28913), .A2(n31208), .B1(n28069), .B2(img[1073]), .O(
        n27150) );
  ND3S U29130 ( .I1(n27156), .I2(n27150), .I3(n27149), .O(n27151) );
  MUX2 U29131 ( .A(img[1097]), .B(n27151), .S(n28768), .O(n12435) );
  AOI22S U29132 ( .A1(n13778), .A2(img[1137]), .B1(n29457), .B2(n31209), .O(
        n27152) );
  ND2S U29133 ( .I1(n27070), .I2(n27152), .O(n27153) );
  AOI22S U29134 ( .A1(n25591), .A2(n31210), .B1(n24313), .B2(img[1033]), .O(
        n27155) );
  ND3S U29135 ( .I1(n27156), .I2(n27155), .I3(n27154), .O(n27157) );
  MUX2 U29136 ( .A(img[1137]), .B(n27157), .S(n28761), .O(n12389) );
  AOI22S U29137 ( .A1(n13778), .A2(img[1009]), .B1(n29096), .B2(n31211), .O(
        n27158) );
  ND2S U29138 ( .I1(n27156), .I2(n27158), .O(n27159) );
  MUX2 U29139 ( .A(img[905]), .B(n27159), .S(n29300), .O(n12621) );
  AOI22S U29140 ( .A1(n24415), .A2(img[905]), .B1(n25591), .B2(n31212), .O(
        n27160) );
  ND2S U29141 ( .I1(n27156), .I2(n27160), .O(n27161) );
  AOI22S U29142 ( .A1(n28442), .A2(img[585]), .B1(n25468), .B2(n31213), .O(
        n27162) );
  ND2S U29143 ( .I1(n27156), .I2(n27162), .O(n27163) );
  MUX2 U29144 ( .A(n27163), .B(img[561]), .S(n28578), .O(n12965) );
  AOI22S U29145 ( .A1(n26822), .A2(img[561]), .B1(n29397), .B2(n31214), .O(
        n27164) );
  ND2S U29146 ( .I1(n27070), .I2(n27164), .O(n27165) );
  MUX2 U29147 ( .A(n27165), .B(img[585]), .S(n28581), .O(n12947) );
  AOI22S U29148 ( .A1(n28347), .A2(img[73]), .B1(n27511), .B2(n31215), .O(
        n27166) );
  ND2S U29149 ( .I1(n27156), .I2(n27166), .O(n27167) );
  MUX2 U29150 ( .A(img[49]), .B(n27167), .S(n28584), .O(n13482) );
  AOI22S U29151 ( .A1(n29072), .A2(img[49]), .B1(n27735), .B2(n31216), .O(
        n27168) );
  ND2S U29152 ( .I1(n27070), .I2(n27168), .O(n27169) );
  AOI22S U29153 ( .A1(n28840), .A2(img[969]), .B1(n27735), .B2(n31217), .O(
        n27171) );
  ND2S U29154 ( .I1(n27156), .I2(n27171), .O(n27172) );
  AOI22S U29155 ( .A1(n26855), .A2(img[945]), .B1(n27735), .B2(n31218), .O(
        n27173) );
  ND2S U29156 ( .I1(n27156), .I2(n27173), .O(n27174) );
  MUX2 U29157 ( .A(img[969]), .B(n27174), .S(n28623), .O(n12557) );
  AOI22S U29158 ( .A1(n27990), .A2(img[201]), .B1(n27735), .B2(n31219), .O(
        n27175) );
  ND2S U29159 ( .I1(n27156), .I2(n27175), .O(n27176) );
  MUX2 U29160 ( .A(img[177]), .B(n27176), .S(n28626), .O(n13355) );
  AOI22S U29161 ( .A1(n13780), .A2(img[177]), .B1(n27735), .B2(n31220), .O(
        n27177) );
  ND2S U29162 ( .I1(n27156), .I2(n27177), .O(n27178) );
  MUX2 U29163 ( .A(img[201]), .B(n27178), .S(n28629), .O(n13325) );
  AOI22S U29164 ( .A1(n28840), .A2(img[329]), .B1(n28862), .B2(n31221), .O(
        n27179) );
  ND2S U29165 ( .I1(n27156), .I2(n27179), .O(n27180) );
  MUX2 U29166 ( .A(img[305]), .B(n27180), .S(n28632), .O(n13221) );
  AOI22S U29167 ( .A1(n26970), .A2(img[305]), .B1(n27735), .B2(n31222), .O(
        n27181) );
  ND2S U29168 ( .I1(n27156), .I2(n27181), .O(n27182) );
  AOI22S U29169 ( .A1(n13776), .A2(img[457]), .B1(n29194), .B2(n31223), .O(
        n27183) );
  ND2S U29170 ( .I1(n27156), .I2(n27183), .O(n27184) );
  AOI22S U29171 ( .A1(n28083), .A2(img[433]), .B1(n23918), .B2(n31224), .O(
        n27185) );
  ND2S U29172 ( .I1(n27156), .I2(n27185), .O(n27186) );
  MUX2 U29173 ( .A(n27186), .B(img[457]), .S(n28641), .O(n13069) );
  AOI22S U29174 ( .A1(n13778), .A2(img[841]), .B1(n13781), .B2(n31225), .O(
        n27187) );
  ND2S U29175 ( .I1(n27156), .I2(n27187), .O(n27188) );
  AOI22S U29176 ( .A1(n13777), .A2(img[817]), .B1(n13781), .B2(n31226), .O(
        n27189) );
  ND2S U29177 ( .I1(n27156), .I2(n27189), .O(n27190) );
  AOI22S U29178 ( .A1(n13771), .A2(img[713]), .B1(n25377), .B2(n31227), .O(
        n27191) );
  ND2S U29179 ( .I1(n27156), .I2(n27191), .O(n27192) );
  AOI22S U29180 ( .A1(n13772), .A2(img[689]), .B1(n28862), .B2(n31228), .O(
        n27193) );
  ND2S U29181 ( .I1(n27156), .I2(n27193), .O(n27194) );
  AOI22S U29182 ( .A1(n13780), .A2(img[569]), .B1(n28862), .B2(n31229), .O(
        n27195) );
  ND2S U29183 ( .I1(n27070), .I2(n27195), .O(n27196) );
  MUX2 U29184 ( .A(n27196), .B(img[577]), .S(n28799), .O(n12949) );
  AOI22S U29185 ( .A1(n27065), .A2(img[577]), .B1(n13781), .B2(n31230), .O(
        n27197) );
  ND2S U29186 ( .I1(n27156), .I2(n27197), .O(n27198) );
  MUX2 U29187 ( .A(n27198), .B(img[569]), .S(n29532), .O(n12963) );
  AOI22S U29188 ( .A1(n24415), .A2(img[57]), .B1(n25377), .B2(n31231), .O(
        n27199) );
  ND2S U29189 ( .I1(n27156), .I2(n27199), .O(n27200) );
  MUX2 U29190 ( .A(img[65]), .B(n27200), .S(n28804), .O(n13461) );
  AOI22S U29191 ( .A1(n13773), .A2(img[65]), .B1(n29530), .B2(n31232), .O(
        n27201) );
  ND2S U29192 ( .I1(n27156), .I2(n27201), .O(n27202) );
  AOI22S U29193 ( .A1(n28083), .A2(img[953]), .B1(n24755), .B2(n31233), .O(
        n27203) );
  ND2S U29194 ( .I1(n27156), .I2(n27203), .O(n27204) );
  AOI22S U29195 ( .A1(n27987), .A2(img[961]), .B1(n28182), .B2(n31234), .O(
        n27205) );
  ND2S U29196 ( .I1(n27156), .I2(n27205), .O(n27206) );
  MUX2 U29197 ( .A(img[953]), .B(n27206), .S(n28842), .O(n12573) );
  AOI22S U29198 ( .A1(n26855), .A2(img[185]), .B1(n28938), .B2(n31235), .O(
        n27207) );
  ND2S U29199 ( .I1(n27156), .I2(n27207), .O(n27208) );
  MUX2 U29200 ( .A(img[193]), .B(n27208), .S(n28845), .O(n13339) );
  AOI22S U29201 ( .A1(n29435), .A2(img[193]), .B1(n28862), .B2(n31236), .O(
        n27209) );
  ND2S U29202 ( .I1(n27156), .I2(n27209), .O(n27210) );
  MUX2 U29203 ( .A(img[185]), .B(n27210), .S(n28848), .O(n13341) );
  AOI22S U29204 ( .A1(n13772), .A2(img[313]), .B1(n25591), .B2(n31237), .O(
        n27211) );
  ND2S U29205 ( .I1(n27156), .I2(n27211), .O(n27212) );
  MUX2 U29206 ( .A(img[321]), .B(n27212), .S(n28851), .O(n13205) );
  AOI22S U29207 ( .A1(n28442), .A2(img[321]), .B1(n24374), .B2(n31238), .O(
        n27213) );
  ND2S U29208 ( .I1(n27156), .I2(n27213), .O(n27214) );
  AOI22S U29209 ( .A1(n28442), .A2(img[441]), .B1(n25377), .B2(n31239), .O(
        n27215) );
  ND2S U29210 ( .I1(n27156), .I2(n27215), .O(n27216) );
  MUX2 U29211 ( .A(img[449]), .B(n27216), .S(n28857), .O(n13083) );
  AOI22S U29212 ( .A1(n28106), .A2(img[449]), .B1(n29457), .B2(n31240), .O(
        n27217) );
  ND2S U29213 ( .I1(n27156), .I2(n27217), .O(n27218) );
  INV1S U29214 ( .I(img[833]), .O(n27219) );
  AOI22S U29215 ( .A1(n25595), .A2(img[825]), .B1(n28862), .B2(n27219), .O(
        n27220) );
  ND2S U29216 ( .I1(n27156), .I2(n27220), .O(n27221) );
  MUX2 U29217 ( .A(n27221), .B(img[833]), .S(n28879), .O(n12693) );
  INV1S U29218 ( .I(img[825]), .O(n27222) );
  AOI22S U29219 ( .A1(n26101), .A2(img[833]), .B1(n28433), .B2(n27222), .O(
        n27223) );
  ND2S U29220 ( .I1(n27156), .I2(n27223), .O(n27224) );
  AOI22S U29221 ( .A1(n28382), .A2(img[697]), .B1(n28433), .B2(n31241), .O(
        n27225) );
  ND2S U29222 ( .I1(n27156), .I2(n27225), .O(n27226) );
  AOI22S U29223 ( .A1(n25810), .A2(img[705]), .B1(n29530), .B2(n31242), .O(
        n27227) );
  ND2S U29224 ( .I1(n27156), .I2(n27227), .O(n27228) );
  AOI22S U29225 ( .A1(n29435), .A2(img[529]), .B1(n29407), .B2(n31243), .O(
        n27229) );
  ND2S U29226 ( .I1(n27156), .I2(n27229), .O(n27230) );
  MUX2 U29227 ( .A(n27230), .B(img[617]), .S(n29024), .O(n12915) );
  AOI22S U29228 ( .A1(n28083), .A2(img[617]), .B1(n25062), .B2(n31244), .O(
        n27231) );
  ND2S U29229 ( .I1(n27070), .I2(n27231), .O(n27232) );
  AOI22S U29230 ( .A1(n13776), .A2(img[17]), .B1(n25859), .B2(n31245), .O(
        n27233) );
  ND2S U29231 ( .I1(n27070), .I2(n27233), .O(n27234) );
  AOI22S U29232 ( .A1(n29435), .A2(img[105]), .B1(n25591), .B2(n31246), .O(
        n27235) );
  ND2S U29233 ( .I1(n27070), .I2(n27235), .O(n27236) );
  MUX2 U29234 ( .A(img[17]), .B(n27236), .S(n29027), .O(n13509) );
  AOI22S U29235 ( .A1(n28347), .A2(img[913]), .B1(n24755), .B2(n31247), .O(
        n27237) );
  ND2S U29236 ( .I1(n27156), .I2(n27237), .O(n27238) );
  AOI22S U29237 ( .A1(n27987), .A2(img[1001]), .B1(n13781), .B2(n31248), .O(
        n27239) );
  ND2S U29238 ( .I1(n27156), .I2(n27239), .O(n27240) );
  MUX2 U29239 ( .A(img[913]), .B(n27240), .S(n29061), .O(n12619) );
  AOI22S U29240 ( .A1(n29414), .A2(img[145]), .B1(n27511), .B2(n31249), .O(
        n27241) );
  ND2S U29241 ( .I1(n27070), .I2(n27241), .O(n27242) );
  MUX2 U29242 ( .A(img[233]), .B(n27242), .S(n29070), .O(n13293) );
  AOI22S U29243 ( .A1(n28347), .A2(img[233]), .B1(n27511), .B2(n31250), .O(
        n27243) );
  ND2S U29244 ( .I1(n27156), .I2(n27243), .O(n27244) );
  MUX2 U29245 ( .A(img[145]), .B(n27244), .S(n29067), .O(n13387) );
  AOI22S U29246 ( .A1(n25810), .A2(img[273]), .B1(n28037), .B2(n31251), .O(
        n27245) );
  ND2S U29247 ( .I1(n27156), .I2(n27245), .O(n27246) );
  MUX2 U29248 ( .A(img[361]), .B(n27246), .S(n29078), .O(n13171) );
  AOI22S U29249 ( .A1(n27990), .A2(img[361]), .B1(n27049), .B2(n31252), .O(
        n27247) );
  ND2S U29250 ( .I1(n27156), .I2(n27247), .O(n27248) );
  AOI22S U29251 ( .A1(n25810), .A2(img[401]), .B1(n13781), .B2(n31253), .O(
        n27249) );
  ND2S U29252 ( .I1(n27156), .I2(n27249), .O(n27250) );
  MUX2 U29253 ( .A(img[489]), .B(n27250), .S(n29084), .O(n13037) );
  AOI22S U29254 ( .A1(n27957), .A2(img[489]), .B1(n13775), .B2(n31254), .O(
        n27251) );
  ND2S U29255 ( .I1(n27156), .I2(n27251), .O(n27252) );
  INV1S U29256 ( .I(img[873]), .O(n27253) );
  AOI22S U29257 ( .A1(n27110), .A2(img[785]), .B1(n25062), .B2(n27253), .O(
        n27254) );
  ND2S U29258 ( .I1(n27156), .I2(n27254), .O(n27255) );
  AOI22S U29259 ( .A1(n25810), .A2(img[873]), .B1(n27511), .B2(n31255), .O(
        n27256) );
  ND2S U29260 ( .I1(n27070), .I2(n27256), .O(n27257) );
  MUX2 U29261 ( .A(img[785]), .B(n27257), .S(n29102), .O(n12741) );
  AOI22S U29262 ( .A1(n27722), .A2(img[657]), .B1(n29242), .B2(n31256), .O(
        n27258) );
  ND2S U29263 ( .I1(n27070), .I2(n27258), .O(n27259) );
  AOI22S U29264 ( .A1(n27722), .A2(img[745]), .B1(n28592), .B2(n31257), .O(
        n27260) );
  ND2S U29265 ( .I1(n27156), .I2(n27260), .O(n27261) );
  OAI22S U29266 ( .A1(n27263), .A2(n28530), .B1(n13897), .B2(n27262), .O(
        n27264) );
  ND2S U29267 ( .I1(n28550), .I2(A67_shift[75]), .O(n27268) );
  AOI22S U29268 ( .A1(n28554), .A2(A67_shift[107]), .B1(n28551), .B2(
        A67_shift[203]), .O(n27267) );
  NR2 U29269 ( .I1(n27270), .I2(n27269), .O(n27273) );
  AOI22S U29270 ( .A1(n28546), .A2(A67_shift[171]), .B1(n28545), .B2(
        A67_shift[43]), .O(n27271) );
  ND2S U29271 ( .I1(n28550), .I2(A67_shift[91]), .O(n27275) );
  AOI22S U29272 ( .A1(n28554), .A2(A67_shift[123]), .B1(n28553), .B2(
        A67_shift[27]), .O(n27274) );
  NR2 U29273 ( .I1(n27277), .I2(n27276), .O(n27280) );
  AOI22S U29274 ( .A1(n28546), .A2(A67_shift[187]), .B1(n28545), .B2(
        A67_shift[59]), .O(n27278) );
  ND2S U29275 ( .I1(n28564), .I2(gray_avg_out[3]), .O(n27285) );
  ND2S U29276 ( .I1(n28565), .I2(gray_weight_out[3]), .O(n27284) );
  ND2S U29277 ( .I1(n28566), .I2(gray_max_out[3]), .O(n27283) );
  AOI22S U29278 ( .A1(n25595), .A2(img[531]), .B1(n13775), .B2(n31258), .O(
        n27290) );
  ND2S U29279 ( .I1(n27886), .I2(n27290), .O(n27291) );
  MUX2 U29280 ( .A(n27291), .B(img[619]), .S(n29024), .O(n12913) );
  AOI22S U29281 ( .A1(n26101), .A2(img[619]), .B1(n13775), .B2(n31259), .O(
        n27292) );
  ND2S U29282 ( .I1(n27886), .I2(n27292), .O(n27293) );
  AOI22S U29283 ( .A1(n13771), .A2(img[19]), .B1(n13775), .B2(n31260), .O(
        n27294) );
  ND2S U29284 ( .I1(n13768), .I2(n27294), .O(n27295) );
  MUX2 U29285 ( .A(img[107]), .B(n27295), .S(n29030), .O(n13425) );
  AOI22S U29286 ( .A1(n13771), .A2(img[107]), .B1(n13775), .B2(n31261), .O(
        n27296) );
  ND2S U29287 ( .I1(n27886), .I2(n27296), .O(n27297) );
  AOI22S U29288 ( .A1(n13777), .A2(img[1235]), .B1(n13775), .B2(n31262), .O(
        n27298) );
  ND2S U29289 ( .I1(n13768), .I2(n27298), .O(n27299) );
  MUX2 U29290 ( .A(img[1195]), .B(n27299), .S(n29033), .O(n12335) );
  BUF12CK U29291 ( .I(n27769), .O(n27886) );
  AOI22S U29292 ( .A1(n28913), .A2(n31263), .B1(n24313), .B2(img[1195]), .O(
        n27301) );
  ND3S U29293 ( .I1(n27886), .I2(n27301), .I3(n27300), .O(n27302) );
  MUX2 U29294 ( .A(img[1235]), .B(n27302), .S(n29037), .O(n12297) );
  AOI22S U29295 ( .A1(n28913), .A2(n31264), .B1(n25444), .B2(img[1171]), .O(
        n27304) );
  ND3S U29296 ( .I1(n27886), .I2(n27304), .I3(n27303), .O(n27305) );
  MUX2 U29297 ( .A(img[1259]), .B(n27305), .S(n29044), .O(n12271) );
  AOI22S U29298 ( .A1(n13777), .A2(img[1259]), .B1(n29397), .B2(n31265), .O(
        n27306) );
  ND2S U29299 ( .I1(n27886), .I2(n27306), .O(n27307) );
  AOI22S U29300 ( .A1(n25810), .A2(img[1363]), .B1(n28614), .B2(n31266), .O(
        n27308) );
  ND2S U29301 ( .I1(n27886), .I2(n27308), .O(n27309) );
  MUX2 U29302 ( .A(n27309), .B(img[1323]), .S(n29047), .O(n12209) );
  AOI22S U29303 ( .A1(n28913), .A2(n31267), .B1(n24313), .B2(img[1323]), .O(
        n27311) );
  ND3S U29304 ( .I1(n27886), .I2(n27311), .I3(n27310), .O(n27312) );
  MUX2 U29305 ( .A(img[1363]), .B(n27312), .S(n29051), .O(n12167) );
  AOI22S U29306 ( .A1(n28913), .A2(n31268), .B1(n28069), .B2(img[1299]), .O(
        n27314) );
  ND3S U29307 ( .I1(n27886), .I2(n27314), .I3(n27313), .O(n27315) );
  MUX2 U29308 ( .A(img[1387]), .B(n27315), .S(n29058), .O(n12145) );
  AOI22S U29309 ( .A1(n25595), .A2(img[1387]), .B1(n13781), .B2(n31269), .O(
        n27316) );
  ND2S U29310 ( .I1(n27886), .I2(n27316), .O(n27317) );
  MUX2 U29311 ( .A(n27317), .B(img[1299]), .S(n29054), .O(n12231) );
  AOI22S U29312 ( .A1(n25810), .A2(img[915]), .B1(n29096), .B2(n31270), .O(
        n27318) );
  ND2S U29313 ( .I1(n27886), .I2(n27318), .O(n27319) );
  AOI22S U29314 ( .A1(n25810), .A2(img[1003]), .B1(n25062), .B2(n31271), .O(
        n27320) );
  ND2S U29315 ( .I1(n27886), .I2(n27320), .O(n27321) );
  AOI22S U29316 ( .A1(n25810), .A2(img[147]), .B1(n28862), .B2(n31272), .O(
        n27322) );
  ND2S U29317 ( .I1(n27886), .I2(n27322), .O(n27323) );
  MUX2 U29318 ( .A(img[235]), .B(n27323), .S(n29070), .O(n13295) );
  AOI22S U29319 ( .A1(n28106), .A2(img[235]), .B1(n29397), .B2(n31273), .O(
        n27324) );
  ND2S U29320 ( .I1(n27886), .I2(n27324), .O(n27325) );
  MUX2 U29321 ( .A(img[147]), .B(n27325), .S(n29067), .O(n13385) );
  AOI22S U29322 ( .A1(n28083), .A2(img[275]), .B1(n13775), .B2(n31274), .O(
        n27326) );
  ND2S U29323 ( .I1(n27886), .I2(n27326), .O(n27327) );
  MUX2 U29324 ( .A(img[363]), .B(n27327), .S(n29078), .O(n13169) );
  AOI22S U29325 ( .A1(n28347), .A2(img[363]), .B1(n28162), .B2(n31275), .O(
        n27328) );
  ND2S U29326 ( .I1(n27886), .I2(n27328), .O(n27329) );
  AOI22S U29327 ( .A1(n28347), .A2(img[403]), .B1(n24193), .B2(n31276), .O(
        n27330) );
  ND2S U29328 ( .I1(n27886), .I2(n27330), .O(n27331) );
  AOI22S U29329 ( .A1(n28442), .A2(img[491]), .B1(n25591), .B2(n31277), .O(
        n27332) );
  ND2S U29330 ( .I1(n27886), .I2(n27332), .O(n27333) );
  AOI22S U29331 ( .A1(n28840), .A2(img[1491]), .B1(n28433), .B2(n31278), .O(
        n27334) );
  ND2S U29332 ( .I1(n27886), .I2(n27334), .O(n27335) );
  MUX2 U29333 ( .A(n27335), .B(img[1451]), .S(n29087), .O(n12079) );
  AOI22S U29334 ( .A1(n13779), .A2(n27336), .B1(n24946), .B2(img[1451]), .O(
        n27338) );
  ND3S U29335 ( .I1(n27886), .I2(n27338), .I3(n27337), .O(n27339) );
  MUX2 U29336 ( .A(n27339), .B(img[1491]), .S(n29091), .O(n12041) );
  AOI22S U29337 ( .A1(n25377), .A2(n31279), .B1(n28069), .B2(img[1427]), .O(
        n27341) );
  ND3S U29338 ( .I1(n27886), .I2(n27341), .I3(n27340), .O(n27342) );
  MUX2 U29339 ( .A(img[1515]), .B(n27342), .S(n29099), .O(n12015) );
  AOI22S U29340 ( .A1(n13778), .A2(img[1515]), .B1(n29530), .B2(n31280), .O(
        n27343) );
  ND2S U29341 ( .I1(n27886), .I2(n27343), .O(n27344) );
  AOI22S U29342 ( .A1(n13780), .A2(img[787]), .B1(n28037), .B2(n31281), .O(
        n27345) );
  ND2S U29343 ( .I1(n27886), .I2(n27345), .O(n27346) );
  AOI22S U29344 ( .A1(n13778), .A2(img[875]), .B1(n13781), .B2(n31282), .O(
        n27347) );
  ND2S U29345 ( .I1(n27886), .I2(n27347), .O(n27348) );
  MUX2 U29346 ( .A(img[787]), .B(n27348), .S(n29102), .O(n12743) );
  AOI22S U29347 ( .A1(n13772), .A2(img[659]), .B1(n29530), .B2(n31283), .O(
        n27349) );
  ND2S U29348 ( .I1(n27886), .I2(n27349), .O(n27350) );
  AOI22S U29349 ( .A1(n13780), .A2(img[747]), .B1(n29530), .B2(n31284), .O(
        n27351) );
  ND2S U29350 ( .I1(n27886), .I2(n27351), .O(n27352) );
  AOI22S U29351 ( .A1(n28840), .A2(img[1867]), .B1(n28913), .B2(n31285), .O(
        n27353) );
  ND2S U29352 ( .I1(n27886), .I2(n27353), .O(n27354) );
  MUX2 U29353 ( .A(n27354), .B(img[1843]), .S(n28693), .O(n11687) );
  AOI22S U29354 ( .A1(n25591), .A2(n27355), .B1(n28069), .B2(img[1843]), .O(
        n27357) );
  ND3S U29355 ( .I1(n27886), .I2(n27357), .I3(n27356), .O(n27358) );
  MUX2 U29356 ( .A(img[1867]), .B(n27358), .S(n28698), .O(n11665) );
  AOI22S U29357 ( .A1(n13776), .A2(img[1907]), .B1(n29457), .B2(n31286), .O(
        n27359) );
  ND2S U29358 ( .I1(n27886), .I2(n27359), .O(n27360) );
  MUX2 U29359 ( .A(img[1803]), .B(n27360), .S(n28686), .O(n11729) );
  INV1S U29360 ( .I(img[1907]), .O(n27361) );
  AOI22S U29361 ( .A1(n25591), .A2(n27361), .B1(n25444), .B2(img[1803]), .O(
        n27363) );
  AOI22S U29362 ( .A1(n13905), .A2(img[1867]), .B1(img[1899]), .B2(n13782), 
        .O(n27362) );
  ND3S U29363 ( .I1(n27886), .I2(n27363), .I3(n27362), .O(n27364) );
  AOI22S U29364 ( .A1(n13772), .A2(img[1875]), .B1(n13781), .B2(n31287), .O(
        n27365) );
  ND2S U29365 ( .I1(n27886), .I2(n27365), .O(n27366) );
  MUX2 U29366 ( .A(n27366), .B(img[1835]), .S(n28672), .O(n11697) );
  AOI22S U29367 ( .A1(n25591), .A2(n31288), .B1(n24313), .B2(img[1835]), .O(
        n27368) );
  ND2S U29368 ( .I1(n13770), .I2(img[1899]), .O(n27367) );
  ND3S U29369 ( .I1(n27886), .I2(n27368), .I3(n27367), .O(n27369) );
  MUX2 U29370 ( .A(img[1875]), .B(n27369), .S(n28676), .O(n11655) );
  INV1S U29371 ( .I(img[1899]), .O(n27370) );
  AOI22S U29372 ( .A1(n25591), .A2(n27370), .B1(n24313), .B2(img[1811]), .O(
        n27372) );
  AOI22S U29373 ( .A1(n13904), .A2(img[1875]), .B1(img[1907]), .B2(n13782), 
        .O(n27371) );
  ND3S U29374 ( .I1(n27886), .I2(n27372), .I3(n27371), .O(n27373) );
  MUX2 U29375 ( .A(img[1899]), .B(n27373), .S(n28683), .O(n11633) );
  AOI22S U29376 ( .A1(n13772), .A2(img[1899]), .B1(n27511), .B2(n31289), .O(
        n27374) );
  ND2S U29377 ( .I1(n27886), .I2(n27374), .O(n27375) );
  AOI22S U29378 ( .A1(n13772), .A2(img[1739]), .B1(n29096), .B2(n31290), .O(
        n27376) );
  ND2S U29379 ( .I1(n27886), .I2(n27376), .O(n27377) );
  MUX2 U29380 ( .A(n27377), .B(img[1715]), .S(n28722), .O(n11817) );
  AOI22S U29381 ( .A1(n25591), .A2(n27378), .B1(n28254), .B2(img[1715]), .O(
        n27380) );
  ND2S U29382 ( .I1(n13819), .I2(img[1779]), .O(n27379) );
  ND3S U29383 ( .I1(n27886), .I2(n27380), .I3(n27379), .O(n27381) );
  AOI22S U29384 ( .A1(n13772), .A2(img[1779]), .B1(n28343), .B2(n31291), .O(
        n27382) );
  ND2S U29385 ( .I1(n27886), .I2(n27382), .O(n27383) );
  AOI22S U29386 ( .A1(n28614), .A2(n31292), .B1(n24313), .B2(img[1675]), .O(
        n27385) );
  AOI22S U29387 ( .A1(n29124), .A2(img[1739]), .B1(img[1771]), .B2(n13782), 
        .O(n27384) );
  ND3S U29388 ( .I1(n27886), .I2(n27385), .I3(n27384), .O(n27386) );
  MUX2 U29389 ( .A(img[1779]), .B(n27386), .S(n28719), .O(n11753) );
  AOI22S U29390 ( .A1(n28347), .A2(img[1747]), .B1(n13781), .B2(n31293), .O(
        n27387) );
  ND2S U29391 ( .I1(n27886), .I2(n27387), .O(n27388) );
  MUX2 U29392 ( .A(n27388), .B(img[1707]), .S(n28701), .O(n11823) );
  AOI22S U29393 ( .A1(n28614), .A2(n31294), .B1(n28069), .B2(img[1707]), .O(
        n27390) );
  ND3S U29394 ( .I1(n27886), .I2(n27390), .I3(n27389), .O(n27391) );
  MUX2 U29395 ( .A(img[1747]), .B(n27391), .S(n28705), .O(n11785) );
  AOI22S U29396 ( .A1(n28614), .A2(n31295), .B1(n28069), .B2(img[1683]), .O(
        n27393) );
  AOI22S U29397 ( .A1(n13770), .A2(img[1747]), .B1(img[1779]), .B2(n13782), 
        .O(n27392) );
  AOI22S U29398 ( .A1(n29414), .A2(img[1771]), .B1(n25859), .B2(n31296), .O(
        n27395) );
  ND2S U29399 ( .I1(n27886), .I2(n27395), .O(n27396) );
  AOI22S U29400 ( .A1(n28442), .A2(img[1611]), .B1(n28695), .B2(n31297), .O(
        n27397) );
  ND2S U29401 ( .I1(n27886), .I2(n27397), .O(n27398) );
  MUX2 U29402 ( .A(n27398), .B(img[1587]), .S(n28750), .O(n11943) );
  AOI22S U29403 ( .A1(n28182), .A2(n31298), .B1(n28069), .B2(img[1587]), .O(
        n27400) );
  ND3S U29404 ( .I1(n27886), .I2(n27400), .I3(n27399), .O(n27401) );
  MUX2 U29405 ( .A(img[1611]), .B(n27401), .S(n28754), .O(n11921) );
  AOI22S U29406 ( .A1(n29072), .A2(img[1651]), .B1(n13781), .B2(n31299), .O(
        n27402) );
  ND2S U29407 ( .I1(n27886), .I2(n27402), .O(n27403) );
  AOI22S U29408 ( .A1(n28592), .A2(n31300), .B1(n24313), .B2(img[1547]), .O(
        n27405) );
  AOI22S U29409 ( .A1(n13903), .A2(img[1611]), .B1(img[1643]), .B2(n13782), 
        .O(n27404) );
  ND3S U29410 ( .I1(n27886), .I2(n27405), .I3(n27404), .O(n27406) );
  MUX2 U29411 ( .A(img[1651]), .B(n27406), .S(n28747), .O(n11879) );
  AOI22S U29412 ( .A1(n28347), .A2(img[1619]), .B1(n28162), .B2(n31301), .O(
        n27407) );
  ND2S U29413 ( .I1(n27886), .I2(n27407), .O(n27408) );
  MUX2 U29414 ( .A(n27408), .B(img[1579]), .S(n28729), .O(n11953) );
  AOI22S U29415 ( .A1(n28592), .A2(n31302), .B1(n28069), .B2(img[1579]), .O(
        n27410) );
  ND2S U29416 ( .I1(n13905), .I2(img[1643]), .O(n27409) );
  AOI22S U29417 ( .A1(n28592), .A2(n31303), .B1(n28069), .B2(img[1555]), .O(
        n27413) );
  AOI22S U29418 ( .A1(n29124), .A2(img[1619]), .B1(img[1651]), .B2(n13782), 
        .O(n27412) );
  ND3S U29419 ( .I1(n27886), .I2(n27413), .I3(n27412), .O(n27414) );
  MUX2 U29420 ( .A(img[1643]), .B(n27414), .S(n28740), .O(n11889) );
  AOI22S U29421 ( .A1(n28347), .A2(img[1643]), .B1(n28592), .B2(n31304), .O(
        n27415) );
  ND2S U29422 ( .I1(n13768), .I2(n27415), .O(n27416) );
  MUX2 U29423 ( .A(n27416), .B(img[1555]), .S(n28736), .O(n11975) );
  AOI22S U29424 ( .A1(n27990), .A2(img[1107]), .B1(n27735), .B2(n31305), .O(
        n27417) );
  ND2S U29425 ( .I1(n13768), .I2(n27417), .O(n27418) );
  MUX2 U29426 ( .A(n27418), .B(img[1067]), .S(n29115), .O(n12465) );
  AOI22S U29427 ( .A1(n25062), .A2(n31306), .B1(n28069), .B2(img[1067]), .O(
        n27420) );
  ND3S U29428 ( .I1(n27886), .I2(n27420), .I3(n27419), .O(n27421) );
  MUX2 U29429 ( .A(img[1107]), .B(n27421), .S(n29119), .O(n12423) );
  AOI22S U29430 ( .A1(n25062), .A2(n31307), .B1(n24313), .B2(img[1043]), .O(
        n27423) );
  ND3S U29431 ( .I1(n27886), .I2(n27423), .I3(n27422), .O(n27424) );
  MUX2 U29432 ( .A(img[1131]), .B(n27424), .S(n29127), .O(n12401) );
  AOI22S U29433 ( .A1(n28106), .A2(img[1131]), .B1(n25859), .B2(n31308), .O(
        n27425) );
  ND2S U29434 ( .I1(n27886), .I2(n27425), .O(n27426) );
  AOI22S U29435 ( .A1(n25810), .A2(img[1995]), .B1(n29407), .B2(n31309), .O(
        n27427) );
  ND2S U29436 ( .I1(n27886), .I2(n27427), .O(n27428) );
  MUX2 U29437 ( .A(n27428), .B(img[1971]), .S(n28792), .O(n11561) );
  AOI22S U29438 ( .A1(n27735), .A2(n31310), .B1(n24313), .B2(img[1971]), .O(
        n27430) );
  ND3S U29439 ( .I1(n27886), .I2(n27430), .I3(n27429), .O(n27431) );
  MUX2 U29440 ( .A(img[1995]), .B(n27431), .S(n28796), .O(n11535) );
  AOI22S U29441 ( .A1(n24415), .A2(img[2035]), .B1(n29397), .B2(n31311), .O(
        n27432) );
  ND2S U29442 ( .I1(n27886), .I2(n27432), .O(n27433) );
  MUX2 U29443 ( .A(img[1931]), .B(n27433), .S(n28785), .O(n11599) );
  AOI22S U29444 ( .A1(n27443), .A2(n31312), .B1(n28254), .B2(img[1931]), .O(
        n27435) );
  AOI22S U29445 ( .A1(n13903), .A2(img[1995]), .B1(img[2027]), .B2(n28908), 
        .O(n27434) );
  ND3S U29446 ( .I1(n27886), .I2(n27435), .I3(n27434), .O(n27436) );
  MUX2 U29447 ( .A(img[2035]), .B(n27436), .S(n28789), .O(n11497) );
  AOI22S U29448 ( .A1(n26970), .A2(img[2003]), .B1(n13775), .B2(n31313), .O(
        n27437) );
  ND2S U29449 ( .I1(n27886), .I2(n27437), .O(n27438) );
  AOI22S U29450 ( .A1(n27443), .A2(n31314), .B1(n24313), .B2(img[1963]), .O(
        n27440) );
  ND2S U29451 ( .I1(n13903), .I2(img[2027]), .O(n27439) );
  ND3S U29452 ( .I1(n27886), .I2(n27440), .I3(n27439), .O(n27441) );
  MUX2 U29453 ( .A(img[2003]), .B(n27441), .S(n28775), .O(n11529) );
  INV1S U29454 ( .I(img[2027]), .O(n27442) );
  AOI22S U29455 ( .A1(n27443), .A2(n27442), .B1(n27919), .B2(img[1939]), .O(
        n27445) );
  AOI22S U29456 ( .A1(n13905), .A2(img[2003]), .B1(img[2035]), .B2(n13782), 
        .O(n27444) );
  ND3S U29457 ( .I1(n27886), .I2(n27445), .I3(n27444), .O(n27446) );
  AOI22S U29458 ( .A1(n13772), .A2(img[2027]), .B1(n13779), .B2(n31315), .O(
        n27447) );
  ND2S U29459 ( .I1(n27886), .I2(n27447), .O(n27448) );
  MUX2 U29460 ( .A(n27448), .B(img[1939]), .S(n28778), .O(n11593) );
  AOI22S U29461 ( .A1(n13772), .A2(img[555]), .B1(n25591), .B2(n31316), .O(
        n27449) );
  ND2S U29462 ( .I1(n27886), .I2(n27449), .O(n27450) );
  MUX2 U29463 ( .A(n27450), .B(img[595]), .S(n29133), .O(n12935) );
  AOI22S U29464 ( .A1(n13772), .A2(img[595]), .B1(n28862), .B2(n31317), .O(
        n27451) );
  ND2S U29465 ( .I1(n27886), .I2(n27451), .O(n27452) );
  MUX2 U29466 ( .A(n27452), .B(img[555]), .S(n29439), .O(n12977) );
  AOI22S U29467 ( .A1(n13772), .A2(img[43]), .B1(n27511), .B2(n31318), .O(
        n27453) );
  ND2S U29468 ( .I1(n13768), .I2(n27453), .O(n27454) );
  MUX2 U29469 ( .A(img[83]), .B(n27454), .S(n29139), .O(n13447) );
  AOI22S U29470 ( .A1(n13772), .A2(img[83]), .B1(n28695), .B2(n31319), .O(
        n27455) );
  ND2S U29471 ( .I1(n27886), .I2(n27455), .O(n27456) );
  AOI22S U29472 ( .A1(n13772), .A2(img[939]), .B1(n13781), .B2(n31320), .O(
        n27457) );
  ND2S U29473 ( .I1(n27886), .I2(n27457), .O(n27458) );
  AOI22S U29474 ( .A1(n13772), .A2(img[979]), .B1(n29194), .B2(n31321), .O(
        n27459) );
  ND2S U29475 ( .I1(n27886), .I2(n27459), .O(n27460) );
  AOI22S U29476 ( .A1(n28840), .A2(img[171]), .B1(n13781), .B2(n31322), .O(
        n27461) );
  ND2S U29477 ( .I1(n27886), .I2(n27461), .O(n27462) );
  MUX2 U29478 ( .A(img[211]), .B(n27462), .S(n29151), .O(n13321) );
  AOI22S U29479 ( .A1(n28382), .A2(img[211]), .B1(n28592), .B2(n31323), .O(
        n27463) );
  ND2S U29480 ( .I1(n27886), .I2(n27463), .O(n27464) );
  MUX2 U29481 ( .A(img[171]), .B(n27464), .S(n29148), .O(n13359) );
  AOI22S U29482 ( .A1(n29435), .A2(img[299]), .B1(n28592), .B2(n31324), .O(
        n27465) );
  ND2S U29483 ( .I1(n27886), .I2(n27465), .O(n27466) );
  MUX2 U29484 ( .A(img[339]), .B(n27466), .S(n29157), .O(n13191) );
  AOI22S U29485 ( .A1(n29072), .A2(img[339]), .B1(n25062), .B2(n31325), .O(
        n27467) );
  ND2S U29486 ( .I1(n27886), .I2(n27467), .O(n27468) );
  AOI22S U29487 ( .A1(n29435), .A2(img[427]), .B1(n25062), .B2(n31326), .O(
        n27469) );
  ND2S U29488 ( .I1(n27886), .I2(n27469), .O(n27470) );
  AOI22S U29489 ( .A1(n26855), .A2(img[467]), .B1(n25591), .B2(n31327), .O(
        n27471) );
  ND2S U29490 ( .I1(n27886), .I2(n27471), .O(n27472) );
  AOI22S U29491 ( .A1(n29435), .A2(img[811]), .B1(n27735), .B2(n31328), .O(
        n27473) );
  ND2S U29492 ( .I1(n27886), .I2(n27473), .O(n27474) );
  AOI22S U29493 ( .A1(n25595), .A2(img[851]), .B1(n13775), .B2(n31329), .O(
        n27475) );
  ND2S U29494 ( .I1(n27886), .I2(n27475), .O(n27476) );
  MUX2 U29495 ( .A(n27476), .B(img[811]), .S(n29166), .O(n12721) );
  AOI22S U29496 ( .A1(n28347), .A2(img[683]), .B1(n13781), .B2(n31330), .O(
        n27477) );
  ND2S U29497 ( .I1(n27886), .I2(n27477), .O(n27478) );
  AOI22S U29498 ( .A1(n13771), .A2(img[723]), .B1(n24374), .B2(n31331), .O(
        n27479) );
  ND2S U29499 ( .I1(n27886), .I2(n27479), .O(n27480) );
  AOI22S U29500 ( .A1(n28347), .A2(img[579]), .B1(n28695), .B2(n31332), .O(
        n27481) );
  ND2S U29501 ( .I1(n13768), .I2(n27481), .O(n27482) );
  MUX2 U29502 ( .A(n27482), .B(img[571]), .S(n29532), .O(n12961) );
  AOI22S U29503 ( .A1(n13777), .A2(img[571]), .B1(n29397), .B2(n31333), .O(
        n27483) );
  ND2S U29504 ( .I1(n13768), .I2(n27483), .O(n27484) );
  MUX2 U29505 ( .A(n27484), .B(img[579]), .S(n28799), .O(n12951) );
  AOI22S U29506 ( .A1(n13777), .A2(img[67]), .B1(n25591), .B2(n31334), .O(
        n27485) );
  ND2S U29507 ( .I1(n13768), .I2(n27485), .O(n27486) );
  MUX2 U29508 ( .A(img[59]), .B(n27486), .S(n28807), .O(n13473) );
  AOI22S U29509 ( .A1(n13777), .A2(img[59]), .B1(n13781), .B2(n31335), .O(
        n27487) );
  ND2S U29510 ( .I1(n13768), .I2(n27487), .O(n27488) );
  MUX2 U29511 ( .A(img[67]), .B(n27488), .S(n28804), .O(n13463) );
  AOI22S U29512 ( .A1(n13777), .A2(img[1275]), .B1(n28037), .B2(n31336), .O(
        n27489) );
  ND2S U29513 ( .I1(n13768), .I2(n27489), .O(n27490) );
  MUX2 U29514 ( .A(img[1155]), .B(n27490), .S(n28810), .O(n12377) );
  AOI22S U29515 ( .A1(n29194), .A2(n31337), .B1(n28069), .B2(img[1155]), .O(
        n27492) );
  ND3S U29516 ( .I1(n27886), .I2(n27492), .I3(n27491), .O(n27493) );
  MUX2 U29517 ( .A(img[1275]), .B(n27493), .S(n28814), .O(n12255) );
  AOI22S U29518 ( .A1(n27990), .A2(img[1219]), .B1(n28343), .B2(n31338), .O(
        n27494) );
  ND2S U29519 ( .I1(n13768), .I2(n27494), .O(n27495) );
  MUX2 U29520 ( .A(img[1211]), .B(n27495), .S(n28821), .O(n12319) );
  AOI22S U29521 ( .A1(n28135), .A2(n31339), .B1(n28069), .B2(img[1211]), .O(
        n27497) );
  ND3S U29522 ( .I1(n27886), .I2(n27497), .I3(n27496), .O(n27498) );
  MUX2 U29523 ( .A(img[1219]), .B(n27498), .S(n28818), .O(n12313) );
  AOI22S U29524 ( .A1(n29072), .A2(img[1403]), .B1(n29096), .B2(n31340), .O(
        n27499) );
  ND2S U29525 ( .I1(n13768), .I2(n27499), .O(n27500) );
  MUX2 U29526 ( .A(img[1283]), .B(n27500), .S(n28824), .O(n12247) );
  AOI22S U29527 ( .A1(n28592), .A2(n31341), .B1(n28069), .B2(img[1283]), .O(
        n27502) );
  ND3S U29528 ( .I1(n27886), .I2(n27502), .I3(n27501), .O(n27503) );
  MUX2 U29529 ( .A(img[1403]), .B(n27503), .S(n28828), .O(n12129) );
  AOI22S U29530 ( .A1(n27746), .A2(img[1347]), .B1(n27511), .B2(n31342), .O(
        n27504) );
  ND2S U29531 ( .I1(n13768), .I2(n27504), .O(n27505) );
  AOI22S U29532 ( .A1(n28343), .A2(n31343), .B1(n28254), .B2(img[1339]), .O(
        n27507) );
  ND3S U29533 ( .I1(n27886), .I2(n27507), .I3(n27506), .O(n27508) );
  MUX2 U29534 ( .A(img[1347]), .B(n27508), .S(n28832), .O(n12183) );
  AOI22S U29535 ( .A1(n28083), .A2(img[963]), .B1(n27511), .B2(n31344), .O(
        n27509) );
  ND2S U29536 ( .I1(n13768), .I2(n27509), .O(n27510) );
  AOI22S U29537 ( .A1(n13780), .A2(img[955]), .B1(n27511), .B2(n31345), .O(
        n27512) );
  ND2S U29538 ( .I1(n13768), .I2(n27512), .O(n27513) );
  MUX2 U29539 ( .A(img[963]), .B(n27513), .S(n28838), .O(n12569) );
  AOI22S U29540 ( .A1(n29072), .A2(img[195]), .B1(n25062), .B2(n31346), .O(
        n27514) );
  ND2S U29541 ( .I1(n13768), .I2(n27514), .O(n27515) );
  MUX2 U29542 ( .A(img[187]), .B(n27515), .S(n28848), .O(n13343) );
  AOI22S U29543 ( .A1(n29414), .A2(img[187]), .B1(n29407), .B2(n31347), .O(
        n27516) );
  ND2S U29544 ( .I1(n13768), .I2(n27516), .O(n27517) );
  MUX2 U29545 ( .A(img[195]), .B(n27517), .S(n28845), .O(n13337) );
  AOI22S U29546 ( .A1(n28083), .A2(img[323]), .B1(n13781), .B2(n31348), .O(
        n27518) );
  ND2S U29547 ( .I1(n13768), .I2(n27518), .O(n27519) );
  AOI22S U29548 ( .A1(n13776), .A2(img[315]), .B1(n25859), .B2(n31349), .O(
        n27520) );
  ND2S U29549 ( .I1(n13768), .I2(n27520), .O(n27521) );
  MUX2 U29550 ( .A(img[323]), .B(n27521), .S(n28851), .O(n13207) );
  AOI22S U29551 ( .A1(n13771), .A2(img[451]), .B1(n24374), .B2(n31350), .O(
        n27522) );
  ND2S U29552 ( .I1(n13768), .I2(n27522), .O(n27523) );
  MUX2 U29553 ( .A(img[443]), .B(n27523), .S(n28860), .O(n13088) );
  AOI22S U29554 ( .A1(n28442), .A2(img[443]), .B1(n13781), .B2(n31351), .O(
        n27524) );
  ND2S U29555 ( .I1(n13768), .I2(n27524), .O(n27525) );
  MUX2 U29556 ( .A(img[451]), .B(n27525), .S(n28857), .O(n13081) );
  AOI22S U29557 ( .A1(n13777), .A2(img[1531]), .B1(n29096), .B2(n31352), .O(
        n27526) );
  ND2S U29558 ( .I1(n13768), .I2(n27526), .O(n27527) );
  AOI22S U29559 ( .A1(n25062), .A2(n31353), .B1(n28254), .B2(img[1411]), .O(
        n27529) );
  ND3S U29560 ( .I1(n27886), .I2(n27529), .I3(n27528), .O(n27530) );
  MUX2 U29561 ( .A(img[1531]), .B(n27530), .S(n28868), .O(n11999) );
  AOI22S U29562 ( .A1(n13777), .A2(img[1475]), .B1(n25377), .B2(n31354), .O(
        n27531) );
  ND2S U29563 ( .I1(n13768), .I2(n27531), .O(n27532) );
  MUX2 U29564 ( .A(img[1467]), .B(n27532), .S(n28875), .O(n12063) );
  AOI22S U29565 ( .A1(n28343), .A2(n31355), .B1(n28254), .B2(img[1467]), .O(
        n27534) );
  ND3S U29566 ( .I1(n27886), .I2(n27534), .I3(n27533), .O(n27535) );
  MUX2 U29567 ( .A(img[1475]), .B(n27535), .S(n28872), .O(n12057) );
  INV1S U29568 ( .I(img[827]), .O(n27536) );
  AOI22S U29569 ( .A1(n13777), .A2(img[835]), .B1(n28938), .B2(n27536), .O(
        n27537) );
  ND2S U29570 ( .I1(n13768), .I2(n27537), .O(n27538) );
  INV1S U29571 ( .I(img[835]), .O(n27539) );
  AOI22S U29572 ( .A1(n13777), .A2(img[827]), .B1(n28037), .B2(n27539), .O(
        n27540) );
  ND2S U29573 ( .I1(n13768), .I2(n27540), .O(n27541) );
  MUX2 U29574 ( .A(n27541), .B(img[835]), .S(n28879), .O(n12695) );
  AOI22S U29575 ( .A1(n13777), .A2(img[707]), .B1(n28343), .B2(n31356), .O(
        n27542) );
  ND2S U29576 ( .I1(n13768), .I2(n27542), .O(n27543) );
  AOI22S U29577 ( .A1(n13777), .A2(img[699]), .B1(n28433), .B2(n31357), .O(
        n27544) );
  ND2S U29578 ( .I1(n13768), .I2(n27544), .O(n27545) );
  AOI22S U29579 ( .A1(n13777), .A2(img[1883]), .B1(n24193), .B2(n31358), .O(
        n27546) );
  ND2S U29580 ( .I1(n13768), .I2(n27546), .O(n27547) );
  MUX2 U29581 ( .A(n27547), .B(img[1827]), .S(n28892), .O(n11703) );
  AOI22S U29582 ( .A1(n25062), .A2(n31359), .B1(n28069), .B2(img[1827]), .O(
        n27549) );
  ND2S U29583 ( .I1(n29124), .I2(img[1891]), .O(n27548) );
  ND3S U29584 ( .I1(n27886), .I2(n27549), .I3(n27548), .O(n27550) );
  AOI22S U29585 ( .A1(n29435), .A2(img[1891]), .B1(n28433), .B2(n31360), .O(
        n27551) );
  ND2S U29586 ( .I1(n13768), .I2(n27551), .O(n27552) );
  MUX2 U29587 ( .A(img[1819]), .B(n27552), .S(n28899), .O(n11713) );
  AOI22S U29588 ( .A1(n28075), .A2(n31361), .B1(n28069), .B2(img[1819]), .O(
        n27554) );
  AOI22S U29589 ( .A1(n13905), .A2(img[1883]), .B1(img[1915]), .B2(n13782), 
        .O(n27553) );
  ND3S U29590 ( .I1(n27886), .I2(n27554), .I3(n27553), .O(n27555) );
  MUX2 U29591 ( .A(img[1891]), .B(n27555), .S(n28903), .O(n11639) );
  AOI22S U29592 ( .A1(n24415), .A2(img[1915]), .B1(n13781), .B2(n31362), .O(
        n27556) );
  ND2S U29593 ( .I1(n13768), .I2(n27556), .O(n27557) );
  AOI22S U29594 ( .A1(n28913), .A2(n31363), .B1(n28069), .B2(img[1795]), .O(
        n27559) );
  AOI22S U29595 ( .A1(n13905), .A2(img[1859]), .B1(img[1891]), .B2(n13782), 
        .O(n27558) );
  ND3S U29596 ( .I1(n27886), .I2(n27559), .I3(n27558), .O(n27560) );
  MUX2 U29597 ( .A(img[1915]), .B(n27560), .S(n28911), .O(n11617) );
  AOI22S U29598 ( .A1(n26101), .A2(img[1859]), .B1(n28862), .B2(n31364), .O(
        n27561) );
  ND2S U29599 ( .I1(n13768), .I2(n27561), .O(n27562) );
  MUX2 U29600 ( .A(img[1851]), .B(n27562), .S(n28919), .O(n11681) );
  AOI22S U29601 ( .A1(n28343), .A2(n31365), .B1(n24313), .B2(img[1851]), .O(
        n27564) );
  ND3S U29602 ( .I1(n27886), .I2(n27564), .I3(n27563), .O(n27565) );
  MUX2 U29603 ( .A(img[1859]), .B(n27565), .S(n28916), .O(n11671) );
  AOI22S U29604 ( .A1(n28347), .A2(img[1755]), .B1(n13781), .B2(n31366), .O(
        n27566) );
  ND2S U29605 ( .I1(n13768), .I2(n27566), .O(n27567) );
  MUX2 U29606 ( .A(n27567), .B(img[1699]), .S(n28922), .O(n11833) );
  AOI22S U29607 ( .A1(n28938), .A2(n31367), .B1(n28254), .B2(img[1699]), .O(
        n27569) );
  ND3S U29608 ( .I1(n27886), .I2(n27569), .I3(n27568), .O(n27570) );
  AOI22S U29609 ( .A1(n13773), .A2(img[1763]), .B1(n29397), .B2(n31368), .O(
        n27571) );
  ND2S U29610 ( .I1(n13768), .I2(n27571), .O(n27572) );
  MUX2 U29611 ( .A(img[1691]), .B(n27572), .S(n28929), .O(n11839) );
  AOI22S U29612 ( .A1(n29194), .A2(n31369), .B1(n28069), .B2(img[1691]), .O(
        n27574) );
  AOI22S U29613 ( .A1(n13819), .A2(img[1755]), .B1(img[1787]), .B2(n13782), 
        .O(n27573) );
  ND3S U29614 ( .I1(n27886), .I2(n27574), .I3(n27573), .O(n27575) );
  MUX2 U29615 ( .A(img[1763]), .B(n27575), .S(n28933), .O(n11769) );
  AOI22S U29616 ( .A1(n27065), .A2(img[1787]), .B1(n25062), .B2(n31370), .O(
        n27576) );
  ND2S U29617 ( .I1(n13768), .I2(n27576), .O(n27577) );
  AOI22S U29618 ( .A1(n28862), .A2(n31371), .B1(n28069), .B2(img[1667]), .O(
        n27579) );
  AOI22S U29619 ( .A1(n29124), .A2(img[1731]), .B1(img[1763]), .B2(n13782), 
        .O(n27578) );
  ND3S U29620 ( .I1(n27886), .I2(n27579), .I3(n27578), .O(n27580) );
  MUX2 U29621 ( .A(img[1787]), .B(n27580), .S(n28941), .O(n11743) );
  AOI22S U29622 ( .A1(n28412), .A2(img[1731]), .B1(n13781), .B2(n31372), .O(
        n27581) );
  ND2S U29623 ( .I1(n13768), .I2(n27581), .O(n27582) );
  MUX2 U29624 ( .A(img[1723]), .B(n27582), .S(n28948), .O(n11807) );
  AOI22S U29625 ( .A1(n28938), .A2(n31373), .B1(n24313), .B2(img[1723]), .O(
        n27584) );
  ND3S U29626 ( .I1(n27886), .I2(n27584), .I3(n27583), .O(n27585) );
  MUX2 U29627 ( .A(img[1731]), .B(n27585), .S(n28945), .O(n11801) );
  AOI22S U29628 ( .A1(n28347), .A2(img[1627]), .B1(n28075), .B2(n31374), .O(
        n27586) );
  ND2S U29629 ( .I1(n13768), .I2(n27586), .O(n27587) );
  MUX2 U29630 ( .A(n27587), .B(img[1571]), .S(n28951), .O(n11959) );
  AOI22S U29631 ( .A1(n28695), .A2(n27588), .B1(n24946), .B2(img[1571]), .O(
        n27590) );
  ND3S U29632 ( .I1(n27886), .I2(n27590), .I3(n27589), .O(n27591) );
  AOI22S U29633 ( .A1(n29129), .A2(img[1635]), .B1(n27511), .B2(n31375), .O(
        n27592) );
  ND2S U29634 ( .I1(n13768), .I2(n27592), .O(n27593) );
  MUX2 U29635 ( .A(img[1563]), .B(n27593), .S(n28958), .O(n11969) );
  AOI22S U29636 ( .A1(n28938), .A2(n31376), .B1(n24313), .B2(img[1563]), .O(
        n27595) );
  AOI22S U29637 ( .A1(n13903), .A2(img[1627]), .B1(img[1659]), .B2(n13782), 
        .O(n27594) );
  ND3S U29638 ( .I1(n27886), .I2(n27595), .I3(n27594), .O(n27596) );
  MUX2 U29639 ( .A(img[1635]), .B(n27596), .S(n28962), .O(n11894) );
  AOI22S U29640 ( .A1(n26101), .A2(img[1659]), .B1(n28862), .B2(n31377), .O(
        n27597) );
  ND2S U29641 ( .I1(n13768), .I2(n27597), .O(n27598) );
  AOI22S U29642 ( .A1(n29530), .A2(n31378), .B1(n24313), .B2(img[1539]), .O(
        n27600) );
  AOI22S U29643 ( .A1(n13905), .A2(img[1603]), .B1(img[1635]), .B2(n13782), 
        .O(n27599) );
  ND3S U29644 ( .I1(n27886), .I2(n27600), .I3(n27599), .O(n27601) );
  MUX2 U29645 ( .A(img[1659]), .B(n27601), .S(n28969), .O(n11873) );
  AOI22S U29646 ( .A1(n29435), .A2(img[1603]), .B1(n25377), .B2(n31379), .O(
        n27602) );
  ND2S U29647 ( .I1(n13768), .I2(n27602), .O(n27603) );
  AOI22S U29648 ( .A1(n29096), .A2(n31380), .B1(n28069), .B2(img[1595]), .O(
        n27605) );
  ND2S U29649 ( .I1(n29124), .I2(img[1659]), .O(n27604) );
  ND3S U29650 ( .I1(n27886), .I2(n27605), .I3(n27604), .O(n27606) );
  MUX2 U29651 ( .A(img[1603]), .B(n27606), .S(n28973), .O(n11927) );
  AOI22S U29652 ( .A1(n28442), .A2(img[1147]), .B1(n13781), .B2(n31381), .O(
        n27607) );
  ND2S U29653 ( .I1(n13768), .I2(n27607), .O(n27608) );
  MUX2 U29654 ( .A(img[1027]), .B(n27608), .S(n28979), .O(n12503) );
  AOI22S U29655 ( .A1(n23918), .A2(n27609), .B1(n24313), .B2(img[1027]), .O(
        n27611) );
  ND3S U29656 ( .I1(n27886), .I2(n27611), .I3(n27610), .O(n27612) );
  AOI22S U29657 ( .A1(n13772), .A2(img[1091]), .B1(n27735), .B2(n31382), .O(
        n27613) );
  ND2S U29658 ( .I1(n13768), .I2(n27613), .O(n27614) );
  AOI22S U29659 ( .A1(n28182), .A2(n27615), .B1(n24890), .B2(img[1083]), .O(
        n27617) );
  ND2S U29660 ( .I1(n29124), .I2(img[1147]), .O(n27616) );
  ND3S U29661 ( .I1(n27886), .I2(n27617), .I3(n27616), .O(n27618) );
  MUX2 U29662 ( .A(img[1091]), .B(n27618), .S(n28987), .O(n12441) );
  AOI22S U29663 ( .A1(n28347), .A2(img[2011]), .B1(n29407), .B2(n31383), .O(
        n27619) );
  ND2S U29664 ( .I1(n13768), .I2(n27619), .O(n27620) );
  INV1S U29665 ( .I(img[2011]), .O(n27621) );
  AOI22S U29666 ( .A1(n28182), .A2(n27621), .B1(n28043), .B2(img[1955]), .O(
        n27623) );
  ND2S U29667 ( .I1(n13819), .I2(img[2019]), .O(n27622) );
  ND3S U29668 ( .I1(n27886), .I2(n27623), .I3(n27622), .O(n27624) );
  MUX2 U29669 ( .A(img[2011]), .B(n27624), .S(n28997), .O(n11519) );
  AOI22S U29670 ( .A1(n28083), .A2(img[2019]), .B1(n25468), .B2(n31384), .O(
        n27625) );
  ND2S U29671 ( .I1(n13768), .I2(n27625), .O(n27626) );
  MUX2 U29672 ( .A(img[1947]), .B(n27626), .S(n29000), .O(n11583) );
  INV1S U29673 ( .I(img[2019]), .O(n27627) );
  AOI22S U29674 ( .A1(n23918), .A2(n27627), .B1(n28069), .B2(img[1947]), .O(
        n27629) );
  AOI22S U29675 ( .A1(n13905), .A2(img[2011]), .B1(img[2043]), .B2(n13782), 
        .O(n27628) );
  ND3S U29676 ( .I1(n27886), .I2(n27629), .I3(n27628), .O(n27630) );
  AOI22S U29677 ( .A1(n28412), .A2(img[2043]), .B1(n29397), .B2(n31385), .O(
        n27631) );
  ND2S U29678 ( .I1(n13768), .I2(n27631), .O(n27632) );
  MUX2 U29679 ( .A(img[1923]), .B(n27632), .S(n29007), .O(n11609) );
  AOI22S U29680 ( .A1(n28182), .A2(n31386), .B1(n24946), .B2(img[1923]), .O(
        n27634) );
  AOI22S U29681 ( .A1(n13904), .A2(img[1987]), .B1(img[2019]), .B2(n13782), 
        .O(n27633) );
  ND3S U29682 ( .I1(n27886), .I2(n27634), .I3(n27633), .O(n27635) );
  MUX2 U29683 ( .A(img[2043]), .B(n27635), .S(n29011), .O(n11489) );
  AOI22S U29684 ( .A1(n27065), .A2(img[1987]), .B1(n24374), .B2(n31387), .O(
        n27636) );
  ND2S U29685 ( .I1(n13768), .I2(n27636), .O(n27637) );
  MUX2 U29686 ( .A(img[1979]), .B(n27637), .S(n29018), .O(n11551) );
  AOI22S U29687 ( .A1(n28182), .A2(n31388), .B1(n27919), .B2(img[1979]), .O(
        n27639) );
  ND2S U29688 ( .I1(n29124), .I2(img[2043]), .O(n27638) );
  ND3S U29689 ( .I1(n27886), .I2(n27639), .I3(n27638), .O(n27640) );
  MUX2 U29690 ( .A(img[1987]), .B(n27640), .S(n29015), .O(n11545) );
  AOI22S U29691 ( .A1(n26970), .A2(img[523]), .B1(n28614), .B2(n31389), .O(
        n27641) );
  ND2S U29692 ( .I1(n13768), .I2(n27641), .O(n27642) );
  MUX2 U29693 ( .A(n27642), .B(img[627]), .S(n29292), .O(n12903) );
  AOI22S U29694 ( .A1(n13772), .A2(img[627]), .B1(n28614), .B2(n31390), .O(
        n27643) );
  ND2S U29695 ( .I1(n13768), .I2(n27643), .O(n27644) );
  AOI22S U29696 ( .A1(n28106), .A2(img[11]), .B1(n24193), .B2(n31391), .O(
        n27645) );
  ND2S U29697 ( .I1(n13768), .I2(n27645), .O(n27646) );
  MUX2 U29698 ( .A(img[115]), .B(n27646), .S(n29536), .O(n13415) );
  AOI22S U29699 ( .A1(n24415), .A2(img[115]), .B1(n29242), .B2(n31392), .O(
        n27647) );
  ND2S U29700 ( .I1(n13768), .I2(n27647), .O(n27648) );
  AOI22S U29701 ( .A1(n28347), .A2(img[1227]), .B1(n13781), .B2(n31393), .O(
        n27649) );
  ND2S U29702 ( .I1(n13768), .I2(n27649), .O(n27650) );
  AOI22S U29703 ( .A1(n28162), .A2(n31394), .B1(n28254), .B2(img[1203]), .O(
        n27652) );
  ND2S U29704 ( .I1(n29124), .I2(img[1267]), .O(n27651) );
  ND3S U29705 ( .I1(n27886), .I2(n27652), .I3(n27651), .O(n27653) );
  MUX2 U29706 ( .A(img[1227]), .B(n27653), .S(n28602), .O(n12303) );
  AOI22S U29707 ( .A1(n28162), .A2(n31395), .B1(n25444), .B2(img[1163]), .O(
        n27655) );
  ND2S U29708 ( .I1(n13770), .I2(img[1227]), .O(n27654) );
  ND3S U29709 ( .I1(n27886), .I2(n27655), .I3(n27654), .O(n27656) );
  MUX2 U29710 ( .A(img[1267]), .B(n27656), .S(n28595), .O(n12265) );
  AOI22S U29711 ( .A1(n25810), .A2(img[1267]), .B1(n25591), .B2(n31396), .O(
        n27657) );
  ND2S U29712 ( .I1(n13768), .I2(n27657), .O(n27658) );
  AOI22S U29713 ( .A1(n29414), .A2(img[1355]), .B1(n29242), .B2(n31397), .O(
        n27659) );
  ND2S U29714 ( .I1(n13768), .I2(n27659), .O(n27660) );
  MUX2 U29715 ( .A(n27660), .B(img[1331]), .S(n28612), .O(n12199) );
  AOI22S U29716 ( .A1(n28135), .A2(n31398), .B1(n24313), .B2(img[1331]), .O(
        n27662) );
  ND3S U29717 ( .I1(n27886), .I2(n27662), .I3(n27661), .O(n27663) );
  MUX2 U29718 ( .A(img[1355]), .B(n27663), .S(n28617), .O(n12177) );
  AOI22S U29719 ( .A1(n28135), .A2(n31399), .B1(n24890), .B2(img[1291]), .O(
        n27665) );
  ND3S U29720 ( .I1(n27886), .I2(n27665), .I3(n27664), .O(n27666) );
  MUX2 U29721 ( .A(img[1395]), .B(n27666), .S(n28609), .O(n12135) );
  AOI22S U29722 ( .A1(n28347), .A2(img[1395]), .B1(n28135), .B2(n31400), .O(
        n27667) );
  ND2S U29723 ( .I1(n27886), .I2(n27667), .O(n27668) );
  AOI22S U29724 ( .A1(n28083), .A2(img[907]), .B1(n28592), .B2(n31401), .O(
        n27669) );
  ND2S U29725 ( .I1(n27886), .I2(n27669), .O(n27670) );
  MUX2 U29726 ( .A(img[1011]), .B(n27670), .S(n29303), .O(n12521) );
  AOI22S U29727 ( .A1(n13780), .A2(img[1011]), .B1(n28343), .B2(n31402), .O(
        n27671) );
  ND2S U29728 ( .I1(n27886), .I2(n27671), .O(n27672) );
  AOI22S U29729 ( .A1(n28840), .A2(img[139]), .B1(n28135), .B2(n31403), .O(
        n27673) );
  ND2S U29730 ( .I1(n27886), .I2(n27673), .O(n27674) );
  MUX2 U29731 ( .A(img[243]), .B(n27674), .S(n29309), .O(n13289) );
  AOI22S U29732 ( .A1(n13772), .A2(img[243]), .B1(n27049), .B2(n31404), .O(
        n27675) );
  ND2S U29733 ( .I1(n27886), .I2(n27675), .O(n27676) );
  AOI22S U29734 ( .A1(n13772), .A2(img[267]), .B1(n28075), .B2(n31405), .O(
        n27677) );
  ND2S U29735 ( .I1(n27886), .I2(n27677), .O(n27678) );
  AOI22S U29736 ( .A1(n26970), .A2(img[371]), .B1(n29194), .B2(n31406), .O(
        n27679) );
  ND2S U29737 ( .I1(n27886), .I2(n27679), .O(n27680) );
  MUX2 U29738 ( .A(n27680), .B(img[267]), .S(n29312), .O(n13265) );
  AOI22S U29739 ( .A1(n26970), .A2(img[395]), .B1(n29530), .B2(n31407), .O(
        n27681) );
  ND2S U29740 ( .I1(n27886), .I2(n27681), .O(n27682) );
  AOI22S U29741 ( .A1(n27065), .A2(img[499]), .B1(n23918), .B2(n31408), .O(
        n27683) );
  ND2S U29742 ( .I1(n27886), .I2(n27683), .O(n27684) );
  AOI22S U29743 ( .A1(n27990), .A2(img[1483]), .B1(n23918), .B2(n31409), .O(
        n27686) );
  ND2S U29744 ( .I1(n27886), .I2(n27686), .O(n27687) );
  MUX2 U29745 ( .A(img[1459]), .B(n27687), .S(n28652), .O(n12073) );
  AOI22S U29746 ( .A1(n25377), .A2(n27688), .B1(n27919), .B2(img[1459]), .O(
        n27690) );
  ND3S U29747 ( .I1(n27886), .I2(n27690), .I3(n27689), .O(n27691) );
  AOI22S U29748 ( .A1(n27049), .A2(n31410), .B1(n24313), .B2(img[1419]), .O(
        n27693) );
  ND2S U29749 ( .I1(n13819), .I2(img[1483]), .O(n27692) );
  ND3S U29750 ( .I1(n27886), .I2(n27693), .I3(n27692), .O(n27694) );
  MUX2 U29751 ( .A(img[1523]), .B(n27694), .S(n28649), .O(n12009) );
  AOI22S U29752 ( .A1(n24415), .A2(img[1523]), .B1(n27049), .B2(n31411), .O(
        n27695) );
  ND2S U29753 ( .I1(n27886), .I2(n27695), .O(n27696) );
  MUX2 U29754 ( .A(n27696), .B(img[1419]), .S(n28645), .O(n12111) );
  INV1S U29755 ( .I(img[883]), .O(n27697) );
  AOI22S U29756 ( .A1(n27685), .A2(img[779]), .B1(n29457), .B2(n27697), .O(
        n27698) );
  ND2S U29757 ( .I1(n27886), .I2(n27698), .O(n27699) );
  AOI22S U29758 ( .A1(n13776), .A2(img[883]), .B1(n13779), .B2(n31412), .O(
        n27700) );
  ND2S U29759 ( .I1(n27886), .I2(n27700), .O(n27701) );
  MUX2 U29760 ( .A(img[779]), .B(n27701), .S(n29324), .O(n12753) );
  AOI22S U29761 ( .A1(n13778), .A2(img[651]), .B1(n29530), .B2(n31413), .O(
        n27702) );
  ND2S U29762 ( .I1(n27886), .I2(n27702), .O(n27703) );
  AOI22S U29763 ( .A1(n29129), .A2(img[755]), .B1(n29194), .B2(n31414), .O(
        n27704) );
  ND2S U29764 ( .I1(n27886), .I2(n27704), .O(n27705) );
  AOI22S U29765 ( .A1(n25595), .A2(img[1099]), .B1(n25591), .B2(n31415), .O(
        n27706) );
  ND2S U29766 ( .I1(n13768), .I2(n27706), .O(n27707) );
  MUX2 U29767 ( .A(n27707), .B(img[1075]), .S(n28764), .O(n12455) );
  AOI22S U29768 ( .A1(n28695), .A2(n31416), .B1(n27919), .B2(img[1075]), .O(
        n27709) );
  ND3S U29769 ( .I1(n27886), .I2(n27709), .I3(n27708), .O(n27710) );
  MUX2 U29770 ( .A(img[1099]), .B(n27710), .S(n28768), .O(n12433) );
  AOI22S U29771 ( .A1(n29530), .A2(n31417), .B1(n27919), .B2(img[1035]), .O(
        n27712) );
  ND3S U29772 ( .I1(n27886), .I2(n27712), .I3(n27711), .O(n27713) );
  MUX2 U29773 ( .A(img[1139]), .B(n27713), .S(n28761), .O(n12391) );
  AOI22S U29774 ( .A1(n28106), .A2(img[1139]), .B1(n28695), .B2(n31418), .O(
        n27714) );
  ND2S U29775 ( .I1(n27886), .I2(n27714), .O(n27715) );
  AOI22S U29776 ( .A1(n26970), .A2(img[75]), .B1(n28075), .B2(n31419), .O(
        n27716) );
  ND2S U29777 ( .I1(n27886), .I2(n27716), .O(n27717) );
  AOI22S U29778 ( .A1(n29414), .A2(img[51]), .B1(n28135), .B2(n31420), .O(
        n27718) );
  ND2S U29779 ( .I1(n13768), .I2(n27718), .O(n27719) );
  MUX2 U29780 ( .A(img[75]), .B(n27719), .S(n28587), .O(n13457) );
  AOI22S U29781 ( .A1(n26101), .A2(img[971]), .B1(n29242), .B2(n31421), .O(
        n27720) );
  ND2S U29782 ( .I1(n13768), .I2(n27720), .O(n27721) );
  AOI22S U29783 ( .A1(n27685), .A2(img[947]), .B1(n27049), .B2(n31422), .O(
        n27723) );
  ND2S U29784 ( .I1(n27886), .I2(n27723), .O(n27724) );
  MUX2 U29785 ( .A(img[971]), .B(n27724), .S(n28623), .O(n12559) );
  AOI22S U29786 ( .A1(n28106), .A2(img[203]), .B1(n24755), .B2(n31423), .O(
        n27725) );
  ND2S U29787 ( .I1(n27886), .I2(n27725), .O(n27726) );
  MUX2 U29788 ( .A(img[179]), .B(n27726), .S(n28626), .O(n13353) );
  AOI22S U29789 ( .A1(n26822), .A2(img[179]), .B1(n28862), .B2(n31424), .O(
        n27727) );
  ND2S U29790 ( .I1(n27886), .I2(n27727), .O(n27728) );
  MUX2 U29791 ( .A(img[203]), .B(n27728), .S(n28629), .O(n13327) );
  AOI22S U29792 ( .A1(n27110), .A2(img[331]), .B1(n27735), .B2(n31425), .O(
        n27729) );
  ND2S U29793 ( .I1(n13768), .I2(n27729), .O(n27730) );
  MUX2 U29794 ( .A(img[307]), .B(n27730), .S(n28632), .O(n13223) );
  AOI22S U29795 ( .A1(n27685), .A2(img[307]), .B1(n29457), .B2(n31426), .O(
        n27731) );
  ND2S U29796 ( .I1(n13768), .I2(n27731), .O(n27732) );
  AOI22S U29797 ( .A1(n24415), .A2(img[843]), .B1(n27735), .B2(n31427), .O(
        n27733) );
  ND2S U29798 ( .I1(n27886), .I2(n27733), .O(n27734) );
  AOI22S U29799 ( .A1(n26970), .A2(img[819]), .B1(n27735), .B2(n31428), .O(
        n27736) );
  ND2S U29800 ( .I1(n27886), .I2(n27736), .O(n27737) );
  MUX2 U29801 ( .A(n27737), .B(img[843]), .S(n28663), .O(n12689) );
  AOI22S U29802 ( .A1(n27065), .A2(img[715]), .B1(n28695), .B2(n31429), .O(
        n27738) );
  ND2S U29803 ( .I1(n27886), .I2(n27738), .O(n27739) );
  AOI22S U29804 ( .A1(n28347), .A2(img[691]), .B1(n24193), .B2(n31430), .O(
        n27740) );
  ND2S U29805 ( .I1(n27886), .I2(n27740), .O(n27741) );
  AOI22S U29806 ( .A1(n28347), .A2(img[459]), .B1(n28913), .B2(n31431), .O(
        n27742) );
  ND2S U29807 ( .I1(n13768), .I2(n27742), .O(n27743) );
  AOI22S U29808 ( .A1(n27685), .A2(img[435]), .B1(n29530), .B2(n31432), .O(
        n27744) );
  ND2S U29809 ( .I1(n27886), .I2(n27744), .O(n27745) );
  MUX2 U29810 ( .A(n27745), .B(img[459]), .S(n28641), .O(n13071) );
  AOI22S U29811 ( .A1(n13771), .A2(img[587]), .B1(n28135), .B2(n31433), .O(
        n27747) );
  ND2S U29812 ( .I1(n27886), .I2(n27747), .O(n27748) );
  MUX2 U29813 ( .A(n27748), .B(img[563]), .S(n28578), .O(n12967) );
  AOI22S U29814 ( .A1(n13771), .A2(img[563]), .B1(n28695), .B2(n31434), .O(
        n27749) );
  ND2S U29815 ( .I1(n27886), .I2(n27749), .O(n27750) );
  MUX2 U29816 ( .A(n27750), .B(img[587]), .S(n28581), .O(n12945) );
  AOI22S U29817 ( .A1(n13771), .A2(img[475]), .B1(n23918), .B2(n31435), .O(
        n27751) );
  ND2S U29818 ( .I1(n27886), .I2(n27751), .O(n27752) );
  MUX2 U29819 ( .A(img[419]), .B(n27752), .S(n29367), .O(n13113) );
  AOI22S U29820 ( .A1(n13771), .A2(img[419]), .B1(n29407), .B2(n31436), .O(
        n27753) );
  ND2S U29821 ( .I1(n13768), .I2(n27753), .O(n27754) );
  MUX2 U29822 ( .A(img[475]), .B(n27754), .S(n29364), .O(n13055) );
  AOI22S U29823 ( .A1(n26822), .A2(img[1123]), .B1(n25377), .B2(n31437), .O(
        n27755) );
  ND2S U29824 ( .I1(n27886), .I2(n27755), .O(n27756) );
  AOI22S U29825 ( .A1(n28037), .A2(n31438), .B1(n27919), .B2(img[1051]), .O(
        n27758) );
  ND2S U29826 ( .I1(n13820), .I2(img[1115]), .O(n27757) );
  ND3S U29827 ( .I1(n27886), .I2(n27758), .I3(n27757), .O(n27759) );
  MUX2 U29828 ( .A(img[1123]), .B(n27759), .S(n29198), .O(n12407) );
  AOI22S U29829 ( .A1(n28382), .A2(img[1115]), .B1(n28037), .B2(n31439), .O(
        n27760) );
  ND2S U29830 ( .I1(n13768), .I2(n27760), .O(n27761) );
  MUX2 U29831 ( .A(n27761), .B(img[1059]), .S(n29185), .O(n12471) );
  AOI22S U29832 ( .A1(n28075), .A2(n31440), .B1(n27919), .B2(img[1059]), .O(
        n27763) );
  ND3S U29833 ( .I1(n27886), .I2(n27763), .I3(n27762), .O(n27764) );
  MUX2 U29834 ( .A(img[1115]), .B(n27764), .S(n29189), .O(n12417) );
  AOI22S U29835 ( .A1(n26101), .A2(img[547]), .B1(n29530), .B2(n31441), .O(
        n27765) );
  ND2S U29836 ( .I1(n27886), .I2(n27765), .O(n27766) );
  MUX2 U29837 ( .A(n27766), .B(img[603]), .S(n29478), .O(n12929) );
  AOI22S U29838 ( .A1(n25595), .A2(img[91]), .B1(n24755), .B2(n31442), .O(
        n27767) );
  ND2S U29839 ( .I1(n27886), .I2(n27767), .O(n27768) );
  AOI22S U29840 ( .A1(n27685), .A2(img[35]), .B1(n25377), .B2(n31443), .O(
        n27770) );
  ND2S U29841 ( .I1(n13768), .I2(n27770), .O(n27771) );
  MUX2 U29842 ( .A(img[91]), .B(n27771), .S(n29339), .O(n13441) );
  AOI22S U29843 ( .A1(n27685), .A2(img[1251]), .B1(n28075), .B2(n31444), .O(
        n27772) );
  ND2S U29844 ( .I1(n13768), .I2(n27772), .O(n27773) );
  MUX2 U29845 ( .A(img[1179]), .B(n27773), .S(n29214), .O(n12351) );
  AOI22S U29846 ( .A1(n25062), .A2(n31445), .B1(n27919), .B2(img[1179]), .O(
        n27775) );
  ND3S U29847 ( .I1(n27886), .I2(n27775), .I3(n27774), .O(n27776) );
  MUX2 U29848 ( .A(img[1251]), .B(n27776), .S(n29218), .O(n12281) );
  AOI22S U29849 ( .A1(n27746), .A2(img[1243]), .B1(n29096), .B2(n31446), .O(
        n27777) );
  ND2S U29850 ( .I1(n13768), .I2(n27777), .O(n27778) );
  MUX2 U29851 ( .A(n27778), .B(img[1187]), .S(n29207), .O(n12345) );
  AOI22S U29852 ( .A1(n28135), .A2(n31447), .B1(n27919), .B2(img[1187]), .O(
        n27780) );
  ND2S U29853 ( .I1(n13820), .I2(img[1251]), .O(n27779) );
  ND3S U29854 ( .I1(n27886), .I2(n27780), .I3(n27779), .O(n27781) );
  MUX2 U29855 ( .A(img[1243]), .B(n27781), .S(n29211), .O(n12287) );
  AOI22S U29856 ( .A1(n26822), .A2(img[1379]), .B1(n28938), .B2(n31448), .O(
        n27782) );
  ND2S U29857 ( .I1(n13768), .I2(n27782), .O(n27783) );
  MUX2 U29858 ( .A(img[1307]), .B(n27783), .S(n29240), .O(n12225) );
  AOI22S U29859 ( .A1(n28162), .A2(n31449), .B1(n27919), .B2(img[1307]), .O(
        n27785) );
  ND3S U29860 ( .I1(n27886), .I2(n27785), .I3(n27784), .O(n27786) );
  MUX2 U29861 ( .A(img[1379]), .B(n27786), .S(n29245), .O(n12151) );
  AOI22S U29862 ( .A1(n26822), .A2(img[1371]), .B1(n29194), .B2(n31450), .O(
        n27787) );
  ND2S U29863 ( .I1(n13768), .I2(n27787), .O(n27788) );
  MUX2 U29864 ( .A(n27788), .B(img[1315]), .S(n29233), .O(n12215) );
  AOI22S U29865 ( .A1(n27049), .A2(n31451), .B1(n27919), .B2(img[1315]), .O(
        n27790) );
  ND2S U29866 ( .I1(n13819), .I2(img[1379]), .O(n27789) );
  ND3S U29867 ( .I1(n27886), .I2(n27790), .I3(n27789), .O(n27791) );
  MUX2 U29868 ( .A(img[1371]), .B(n27791), .S(n29237), .O(n12161) );
  AOI22S U29869 ( .A1(n28083), .A2(img[987]), .B1(n28614), .B2(n31452), .O(
        n27792) );
  ND2S U29870 ( .I1(n13768), .I2(n27792), .O(n27793) );
  AOI22S U29871 ( .A1(n25810), .A2(img[931]), .B1(n27735), .B2(n31453), .O(
        n27794) );
  ND2S U29872 ( .I1(n13768), .I2(n27794), .O(n27795) );
  MUX2 U29873 ( .A(img[987]), .B(n27795), .S(n29345), .O(n12543) );
  AOI22S U29874 ( .A1(n13771), .A2(img[219]), .B1(n27735), .B2(n31454), .O(
        n27796) );
  ND2S U29875 ( .I1(n13768), .I2(n27796), .O(n27797) );
  MUX2 U29876 ( .A(img[163]), .B(n27797), .S(n29355), .O(n13369) );
  AOI22S U29877 ( .A1(n13771), .A2(img[163]), .B1(n28343), .B2(n31455), .O(
        n27798) );
  ND2S U29878 ( .I1(n13768), .I2(n27798), .O(n27799) );
  MUX2 U29879 ( .A(img[219]), .B(n27799), .S(n29351), .O(n13311) );
  AOI22S U29880 ( .A1(n13771), .A2(img[1507]), .B1(n29397), .B2(n31456), .O(
        n27800) );
  ND2S U29881 ( .I1(n13768), .I2(n27800), .O(n27801) );
  MUX2 U29882 ( .A(n27801), .B(img[1435]), .S(n29255), .O(n12095) );
  AOI22S U29883 ( .A1(n28913), .A2(n31457), .B1(n27919), .B2(img[1435]), .O(
        n27803) );
  ND3S U29884 ( .I1(n27886), .I2(n27803), .I3(n27802), .O(n27804) );
  AOI22S U29885 ( .A1(n13771), .A2(img[1499]), .B1(n29407), .B2(n31458), .O(
        n27805) );
  ND2S U29886 ( .I1(n13768), .I2(n27805), .O(n27806) );
  AOI22S U29887 ( .A1(n28162), .A2(n31459), .B1(n27919), .B2(img[1443]), .O(
        n27808) );
  ND3S U29888 ( .I1(n27886), .I2(n27808), .I3(n27807), .O(n27809) );
  MUX2 U29889 ( .A(img[1499]), .B(n27809), .S(n29252), .O(n12031) );
  AOI22S U29890 ( .A1(n13771), .A2(img[731]), .B1(n23941), .B2(n31460), .O(
        n27810) );
  ND2S U29891 ( .I1(n13768), .I2(n27810), .O(n27811) );
  AOI22S U29892 ( .A1(n13771), .A2(img[675]), .B1(n25591), .B2(n31461), .O(
        n27812) );
  ND2S U29893 ( .I1(n13768), .I2(n27812), .O(n27813) );
  AOI22S U29894 ( .A1(n13771), .A2(img[347]), .B1(n27735), .B2(n31462), .O(
        n27814) );
  ND2S U29895 ( .I1(n13768), .I2(n27814), .O(n27815) );
  AOI22S U29896 ( .A1(n13776), .A2(img[291]), .B1(n24374), .B2(n31463), .O(
        n27816) );
  ND2S U29897 ( .I1(n13768), .I2(n27816), .O(n27817) );
  MUX2 U29898 ( .A(img[347]), .B(n27817), .S(n29358), .O(n13185) );
  AOI22S U29899 ( .A1(n27746), .A2(img[859]), .B1(n25377), .B2(n31464), .O(
        n27818) );
  ND2S U29900 ( .I1(n13768), .I2(n27818), .O(n27819) );
  MUX2 U29901 ( .A(n27819), .B(img[803]), .S(n29374), .O(n12727) );
  AOI22S U29902 ( .A1(n28412), .A2(img[803]), .B1(n25062), .B2(n31465), .O(
        n27820) );
  ND2S U29903 ( .I1(n13768), .I2(n27820), .O(n27821) );
  AOI22S U29904 ( .A1(n29435), .A2(img[507]), .B1(n23941), .B2(n31466), .O(
        n27822) );
  ND2S U29905 ( .I1(n13768), .I2(n27822), .O(n27823) );
  AOI22S U29906 ( .A1(n26855), .A2(img[387]), .B1(n23941), .B2(n31467), .O(
        n27824) );
  ND2S U29907 ( .I1(n13768), .I2(n27824), .O(n27825) );
  MUX2 U29908 ( .A(n27825), .B(img[507]), .S(n29420), .O(n13023) );
  AOI22S U29909 ( .A1(n29072), .A2(img[635]), .B1(n23918), .B2(n31468), .O(
        n27826) );
  ND2S U29910 ( .I1(n13768), .I2(n27826), .O(n27827) );
  AOI22S U29911 ( .A1(n28106), .A2(img[515]), .B1(n29397), .B2(n31469), .O(
        n27828) );
  ND2S U29912 ( .I1(n13768), .I2(n27828), .O(n27829) );
  MUX2 U29913 ( .A(n27829), .B(img[635]), .S(n29386), .O(n12897) );
  AOI22S U29914 ( .A1(n27746), .A2(img[123]), .B1(n25591), .B2(n31470), .O(
        n27830) );
  ND2S U29915 ( .I1(n13768), .I2(n27830), .O(n27831) );
  AOI22S U29916 ( .A1(n28347), .A2(img[3]), .B1(n13781), .B2(n31471), .O(
        n27832) );
  ND2S U29917 ( .I1(n13768), .I2(n27832), .O(n27833) );
  MUX2 U29918 ( .A(img[123]), .B(n27833), .S(n29392), .O(n13409) );
  AOI22S U29919 ( .A1(n28382), .A2(img[1019]), .B1(n28182), .B2(n31472), .O(
        n27834) );
  ND2S U29920 ( .I1(n13768), .I2(n27834), .O(n27835) );
  AOI22S U29921 ( .A1(n28442), .A2(img[899]), .B1(n28182), .B2(n31473), .O(
        n27836) );
  ND2S U29922 ( .I1(n13768), .I2(n27836), .O(n27837) );
  MUX2 U29923 ( .A(img[1019]), .B(n27837), .S(n29399), .O(n12511) );
  AOI22S U29924 ( .A1(n13777), .A2(img[251]), .B1(n28162), .B2(n31474), .O(
        n27838) );
  ND2S U29925 ( .I1(n13768), .I2(n27838), .O(n27839) );
  MUX2 U29926 ( .A(n27839), .B(img[131]), .S(n29402), .O(n13401) );
  AOI22S U29927 ( .A1(n13777), .A2(img[131]), .B1(n28182), .B2(n31475), .O(
        n27840) );
  ND2S U29928 ( .I1(n27886), .I2(n27840), .O(n27841) );
  MUX2 U29929 ( .A(img[251]), .B(n27841), .S(n29405), .O(n13278) );
  AOI22S U29930 ( .A1(n13777), .A2(img[379]), .B1(n13779), .B2(n31476), .O(
        n27842) );
  ND2S U29931 ( .I1(n27886), .I2(n27842), .O(n27843) );
  AOI22S U29932 ( .A1(n13777), .A2(img[259]), .B1(n28182), .B2(n31477), .O(
        n27844) );
  ND2S U29933 ( .I1(n27886), .I2(n27844), .O(n27845) );
  MUX2 U29934 ( .A(img[379]), .B(n27845), .S(n29412), .O(n13153) );
  AOI22S U29935 ( .A1(n13777), .A2(img[891]), .B1(n28162), .B2(n31478), .O(
        n27846) );
  ND2S U29936 ( .I1(n27886), .I2(n27846), .O(n27847) );
  MUX2 U29937 ( .A(img[771]), .B(n27847), .S(n29423), .O(n12759) );
  INV1S U29938 ( .I(img[891]), .O(n27848) );
  AOI22S U29939 ( .A1(n13777), .A2(img[771]), .B1(n28182), .B2(n27848), .O(
        n27849) );
  ND2S U29940 ( .I1(n27886), .I2(n27849), .O(n27850) );
  AOI22S U29941 ( .A1(n13777), .A2(img[763]), .B1(n28182), .B2(n31479), .O(
        n27851) );
  ND2S U29942 ( .I1(n27886), .I2(n27851), .O(n27852) );
  AOI22S U29943 ( .A1(n13777), .A2(img[643]), .B1(n28162), .B2(n31480), .O(
        n27853) );
  ND2S U29944 ( .I1(n27886), .I2(n27853), .O(n27854) );
  AOI22S U29945 ( .A1(n13777), .A2(img[611]), .B1(n28162), .B2(n31481), .O(
        n27855) );
  ND2S U29946 ( .I1(n27886), .I2(n27855), .O(n27856) );
  AOI22S U29947 ( .A1(n13777), .A2(img[539]), .B1(n29407), .B2(n31482), .O(
        n27857) );
  ND2S U29948 ( .I1(n27886), .I2(n27857), .O(n27858) );
  MUX2 U29949 ( .A(n27858), .B(img[611]), .S(n29286), .O(n12919) );
  AOI22S U29950 ( .A1(n13777), .A2(img[99]), .B1(n29407), .B2(n31483), .O(
        n27859) );
  ND2S U29951 ( .I1(n27886), .I2(n27859), .O(n27860) );
  AOI22S U29952 ( .A1(n27065), .A2(img[27]), .B1(n29407), .B2(n31484), .O(
        n27861) );
  ND2S U29953 ( .I1(n27886), .I2(n27861), .O(n27862) );
  MUX2 U29954 ( .A(img[99]), .B(n27862), .S(n29280), .O(n13431) );
  AOI22S U29955 ( .A1(n29435), .A2(img[995]), .B1(n29407), .B2(n31485), .O(
        n27863) );
  ND2S U29956 ( .I1(n27886), .I2(n27863), .O(n27864) );
  AOI22S U29957 ( .A1(n25595), .A2(img[923]), .B1(n29407), .B2(n31486), .O(
        n27865) );
  ND2S U29958 ( .I1(n27886), .I2(n27865), .O(n27866) );
  MUX2 U29959 ( .A(img[995]), .B(n27866), .S(n29224), .O(n12537) );
  AOI22S U29960 ( .A1(n29435), .A2(img[227]), .B1(n29407), .B2(n31487), .O(
        n27867) );
  ND2S U29961 ( .I1(n13768), .I2(n27867), .O(n27868) );
  MUX2 U29962 ( .A(img[155]), .B(n27868), .S(n29264), .O(n13375) );
  AOI22S U29963 ( .A1(n13773), .A2(img[155]), .B1(n29407), .B2(n31488), .O(
        n27869) );
  ND2S U29964 ( .I1(n27886), .I2(n27869), .O(n27870) );
  MUX2 U29965 ( .A(img[227]), .B(n27870), .S(n29267), .O(n13305) );
  AOI22S U29966 ( .A1(n27065), .A2(img[355]), .B1(n29407), .B2(n31489), .O(
        n27871) );
  ND2S U29967 ( .I1(n27886), .I2(n27871), .O(n27872) );
  MUX2 U29968 ( .A(img[283]), .B(n27872), .S(n29179), .O(n13249) );
  AOI22S U29969 ( .A1(n24415), .A2(img[283]), .B1(n29530), .B2(n31490), .O(
        n27873) );
  ND2S U29970 ( .I1(n27886), .I2(n27873), .O(n27874) );
  AOI22S U29971 ( .A1(n29129), .A2(img[483]), .B1(n29530), .B2(n31491), .O(
        n27875) );
  ND2S U29972 ( .I1(n27886), .I2(n27875), .O(n27876) );
  AOI22S U29973 ( .A1(n28468), .A2(img[411]), .B1(n29530), .B2(n31492), .O(
        n27877) );
  ND2S U29974 ( .I1(n27886), .I2(n27877), .O(n27878) );
  AOI22S U29975 ( .A1(n28412), .A2(img[867]), .B1(n29530), .B2(n31493), .O(
        n27879) );
  ND2S U29976 ( .I1(n27886), .I2(n27879), .O(n27880) );
  MUX2 U29977 ( .A(img[795]), .B(n27880), .S(n29227), .O(n12737) );
  AOI22S U29978 ( .A1(n28347), .A2(img[795]), .B1(n29457), .B2(n31494), .O(
        n27881) );
  ND2S U29979 ( .I1(n27886), .I2(n27881), .O(n27882) );
  AOI22S U29980 ( .A1(n27987), .A2(img[739]), .B1(n29457), .B2(n31495), .O(
        n27883) );
  ND2S U29981 ( .I1(n27886), .I2(n27883), .O(n27884) );
  AOI22S U29982 ( .A1(n27987), .A2(img[667]), .B1(n29397), .B2(n31496), .O(
        n27885) );
  ND2S U29983 ( .I1(n27886), .I2(n27885), .O(n27887) );
  OAI22S U29984 ( .A1(n27889), .A2(n28530), .B1(n13897), .B2(n27888), .O(
        n27890) );
  ND2S U29985 ( .I1(n28547), .I2(A67_shift[248]), .O(n27896) );
  AOI22S U29986 ( .A1(n28552), .A2(A67_shift[152]), .B1(n28551), .B2(
        A67_shift[216]), .O(n27895) );
  ND2S U29987 ( .I1(n28554), .I2(A67_shift[120]), .O(n27894) );
  INV1S U29988 ( .I(A67_shift[56]), .O(n27899) );
  AOI22S U29989 ( .A1(n28553), .A2(A67_shift[24]), .B1(n28546), .B2(
        A67_shift[184]), .O(n27898) );
  AOI12HS U29990 ( .B1(n28550), .B2(A67_shift[88]), .A1(n28555), .O(n27897) );
  OAI112HS U29991 ( .C1(n28544), .C2(n27899), .A1(n27898), .B1(n27897), .O(
        n27908) );
  AOI22S U29992 ( .A1(n28546), .A2(A67_shift[168]), .B1(n28545), .B2(
        A67_shift[40]), .O(n27901) );
  ND2S U29993 ( .I1(n28550), .I2(A67_shift[72]), .O(n27905) );
  AOI22S U29994 ( .A1(n28552), .A2(A67_shift[136]), .B1(n28551), .B2(
        A67_shift[200]), .O(n27904) );
  AOI22S U29995 ( .A1(n28554), .A2(A67_shift[104]), .B1(n28553), .B2(
        A67_shift[8]), .O(n27902) );
  OAI22S U29996 ( .A1(n27909), .A2(n27908), .B1(n27907), .B2(n27906), .O(
        n27914) );
  ND2S U29997 ( .I1(n28564), .I2(gray_avg_out[0]), .O(n27912) );
  ND2S U29998 ( .I1(n28565), .I2(gray_weight_out[0]), .O(n27911) );
  ND2S U29999 ( .I1(n28566), .I2(gray_max_out[0]), .O(n27910) );
  AOI22S U30000 ( .A1(n27987), .A2(img[1272]), .B1(n29407), .B2(n31497), .O(
        n27917) );
  ND2S U30001 ( .I1(n28425), .I2(n27917), .O(n27918) );
  AOI22S U30002 ( .A1(n28162), .A2(n31498), .B1(n27919), .B2(img[1152]), .O(
        n27921) );
  ND3S U30003 ( .I1(n28425), .I2(n27921), .I3(n27920), .O(n27922) );
  MUX2 U30004 ( .A(img[1272]), .B(n27922), .S(n28814), .O(n12260) );
  AOI22S U30005 ( .A1(n27987), .A2(img[1216]), .B1(n29407), .B2(n31499), .O(
        n27923) );
  ND2S U30006 ( .I1(n28425), .I2(n27923), .O(n27924) );
  MUX2 U30007 ( .A(img[1208]), .B(n27924), .S(n28821), .O(n12324) );
  AOI22S U30008 ( .A1(n29242), .A2(n31500), .B1(n27919), .B2(img[1208]), .O(
        n27926) );
  ND3S U30009 ( .I1(n28425), .I2(n27926), .I3(n27925), .O(n27927) );
  MUX2 U30010 ( .A(img[1216]), .B(n27927), .S(n28818), .O(n12316) );
  AOI22S U30011 ( .A1(n13777), .A2(img[1880]), .B1(n29407), .B2(n31501), .O(
        n27928) );
  ND2S U30012 ( .I1(n28425), .I2(n27928), .O(n27929) );
  AOI22S U30013 ( .A1(n27735), .A2(n31502), .B1(n27919), .B2(img[1824]), .O(
        n27931) );
  ND3S U30014 ( .I1(n28425), .I2(n27931), .I3(n27930), .O(n27932) );
  MUX2 U30015 ( .A(img[1880]), .B(n27932), .S(n28896), .O(n11652) );
  AOI22S U30016 ( .A1(n28468), .A2(img[1888]), .B1(n29397), .B2(n31503), .O(
        n27933) );
  ND2S U30017 ( .I1(n28425), .I2(n27933), .O(n27934) );
  AOI22S U30018 ( .A1(n25062), .A2(n31504), .B1(n27919), .B2(img[1816]), .O(
        n27936) );
  AOI22S U30019 ( .A1(n13905), .A2(img[1880]), .B1(img[1912]), .B2(n13782), 
        .O(n27935) );
  ND3S U30020 ( .I1(n28425), .I2(n27936), .I3(n27935), .O(n27937) );
  MUX2 U30021 ( .A(img[1888]), .B(n27937), .S(n28903), .O(n11644) );
  AOI22S U30022 ( .A1(n29435), .A2(img[1912]), .B1(n25591), .B2(n31505), .O(
        n27938) );
  ND2S U30023 ( .I1(n28425), .I2(n27938), .O(n27939) );
  AOI22S U30024 ( .A1(n25591), .A2(n31506), .B1(n27919), .B2(img[1792]), .O(
        n27941) );
  AOI22S U30025 ( .A1(n13905), .A2(img[1856]), .B1(img[1888]), .B2(n13782), 
        .O(n27940) );
  ND3S U30026 ( .I1(n28425), .I2(n27941), .I3(n27940), .O(n27942) );
  MUX2 U30027 ( .A(img[1912]), .B(n27942), .S(n28911), .O(n11620) );
  AOI22S U30028 ( .A1(n28347), .A2(img[1856]), .B1(n25591), .B2(n31507), .O(
        n27943) );
  ND2S U30029 ( .I1(n28425), .I2(n27943), .O(n27944) );
  MUX2 U30030 ( .A(img[1848]), .B(n27944), .S(n28919), .O(n11684) );
  AOI22S U30031 ( .A1(n28862), .A2(n31508), .B1(n27919), .B2(img[1848]), .O(
        n27946) );
  ND3S U30032 ( .I1(n28425), .I2(n27946), .I3(n27945), .O(n27947) );
  MUX2 U30033 ( .A(img[1856]), .B(n27947), .S(n28916), .O(n11676) );
  AOI22S U30034 ( .A1(n13773), .A2(img[576]), .B1(n28913), .B2(n31509), .O(
        n27948) );
  ND2S U30035 ( .I1(n28425), .I2(n27948), .O(n27949) );
  MUX2 U30036 ( .A(n27949), .B(img[568]), .S(n29532), .O(n12964) );
  AOI22S U30037 ( .A1(n26490), .A2(img[568]), .B1(n25591), .B2(n31510), .O(
        n27950) );
  ND2S U30038 ( .I1(n28425), .I2(n27950), .O(n27951) );
  MUX2 U30039 ( .A(n27951), .B(img[576]), .S(n28799), .O(n12956) );
  AOI22S U30040 ( .A1(n29435), .A2(img[1528]), .B1(n28913), .B2(n31511), .O(
        n27952) );
  ND2S U30041 ( .I1(n28425), .I2(n27952), .O(n27953) );
  MUX2 U30042 ( .A(img[1408]), .B(n27953), .S(n28864), .O(n12124) );
  BUF12CK U30043 ( .I(n28415), .O(n28425) );
  AOI22S U30044 ( .A1(n29194), .A2(n31512), .B1(n24313), .B2(img[1408]), .O(
        n27955) );
  ND3S U30045 ( .I1(n28425), .I2(n27955), .I3(n27954), .O(n27956) );
  AOI22S U30046 ( .A1(n26101), .A2(img[1472]), .B1(n28695), .B2(n31513), .O(
        n27958) );
  ND2S U30047 ( .I1(n28425), .I2(n27958), .O(n27959) );
  AOI22S U30048 ( .A1(n29530), .A2(n31514), .B1(n27919), .B2(img[1464]), .O(
        n27961) );
  ND2S U30049 ( .I1(n13770), .I2(img[1528]), .O(n27960) );
  AOI22S U30050 ( .A1(n28347), .A2(img[64]), .B1(n28433), .B2(n31515), .O(
        n27963) );
  ND2S U30051 ( .I1(n28425), .I2(n27963), .O(n27964) );
  AOI22S U30052 ( .A1(n26970), .A2(img[56]), .B1(n27735), .B2(n31516), .O(
        n27965) );
  ND2S U30053 ( .I1(n28425), .I2(n27965), .O(n27966) );
  MUX2 U30054 ( .A(img[64]), .B(n27966), .S(n28804), .O(n13468) );
  AOI22S U30055 ( .A1(n28442), .A2(img[1400]), .B1(n29457), .B2(n31517), .O(
        n27967) );
  ND2S U30056 ( .I1(n28425), .I2(n27967), .O(n27968) );
  MUX2 U30057 ( .A(img[1280]), .B(n27968), .S(n28824), .O(n12252) );
  AOI22S U30058 ( .A1(n28862), .A2(n31518), .B1(n27919), .B2(img[1280]), .O(
        n27970) );
  ND3S U30059 ( .I1(n28425), .I2(n27970), .I3(n27969), .O(n27971) );
  MUX2 U30060 ( .A(img[1400]), .B(n27971), .S(n28828), .O(n12132) );
  AOI22S U30061 ( .A1(n27987), .A2(img[1344]), .B1(n27511), .B2(n31519), .O(
        n27972) );
  ND2S U30062 ( .I1(n28425), .I2(n27972), .O(n27973) );
  AOI22S U30063 ( .A1(n29194), .A2(n31520), .B1(n27919), .B2(img[1336]), .O(
        n27975) );
  ND3S U30064 ( .I1(n28425), .I2(n27975), .I3(n27974), .O(n27976) );
  MUX2 U30065 ( .A(img[1344]), .B(n27976), .S(n28832), .O(n12188) );
  AOI22S U30066 ( .A1(n27987), .A2(img[960]), .B1(n29530), .B2(n31521), .O(
        n27977) );
  ND2S U30067 ( .I1(n28425), .I2(n27977), .O(n27978) );
  MUX2 U30068 ( .A(img[952]), .B(n27978), .S(n28842), .O(n12580) );
  AOI22S U30069 ( .A1(n27987), .A2(img[952]), .B1(n25859), .B2(n31522), .O(
        n27979) );
  ND2S U30070 ( .I1(n28425), .I2(n27979), .O(n27980) );
  AOI22S U30071 ( .A1(n27987), .A2(img[192]), .B1(n28037), .B2(n31523), .O(
        n27981) );
  ND2S U30072 ( .I1(n28425), .I2(n27981), .O(n27982) );
  MUX2 U30073 ( .A(img[184]), .B(n27982), .S(n28848), .O(n13348) );
  AOI22S U30074 ( .A1(n27987), .A2(img[184]), .B1(n23918), .B2(n31524), .O(
        n27983) );
  ND2S U30075 ( .I1(n28425), .I2(n27983), .O(n27984) );
  MUX2 U30076 ( .A(img[192]), .B(n27984), .S(n28845), .O(n13340) );
  AOI22S U30077 ( .A1(n27987), .A2(img[320]), .B1(n25591), .B2(n31525), .O(
        n27985) );
  ND2S U30078 ( .I1(n28425), .I2(n27985), .O(n27986) );
  AOI22S U30079 ( .A1(n27987), .A2(img[312]), .B1(n29407), .B2(n31526), .O(
        n27988) );
  ND2S U30080 ( .I1(n28425), .I2(n27988), .O(n27989) );
  MUX2 U30081 ( .A(img[320]), .B(n27989), .S(n28851), .O(n13212) );
  AOI22S U30082 ( .A1(n13778), .A2(img[448]), .B1(n28862), .B2(n31527), .O(
        n27991) );
  ND2S U30083 ( .I1(n28425), .I2(n27991), .O(n27992) );
  AOI22S U30084 ( .A1(n13778), .A2(img[440]), .B1(n29530), .B2(n31528), .O(
        n27993) );
  ND2S U30085 ( .I1(n28425), .I2(n27993), .O(n27994) );
  INV1S U30086 ( .I(img[824]), .O(n27995) );
  AOI22S U30087 ( .A1(n13778), .A2(img[832]), .B1(n13781), .B2(n27995), .O(
        n27996) );
  ND2S U30088 ( .I1(n28425), .I2(n27996), .O(n27997) );
  INV1S U30089 ( .I(img[832]), .O(n27998) );
  AOI22S U30090 ( .A1(n13778), .A2(img[824]), .B1(n25377), .B2(n27998), .O(
        n27999) );
  ND2S U30091 ( .I1(n28425), .I2(n27999), .O(n28000) );
  MUX2 U30092 ( .A(n28000), .B(img[832]), .S(n28879), .O(n12700) );
  AOI22S U30093 ( .A1(n26101), .A2(img[704]), .B1(n28862), .B2(n31529), .O(
        n28001) );
  ND2S U30094 ( .I1(n28425), .I2(n28001), .O(n28002) );
  AOI22S U30095 ( .A1(n28106), .A2(img[696]), .B1(n25377), .B2(n31530), .O(
        n28003) );
  ND2S U30096 ( .I1(n28425), .I2(n28003), .O(n28004) );
  AOI22S U30097 ( .A1(n25595), .A2(img[1752]), .B1(n28862), .B2(n31531), .O(
        n28005) );
  ND2S U30098 ( .I1(n28425), .I2(n28005), .O(n28006) );
  MUX2 U30099 ( .A(n28006), .B(img[1696]), .S(n28922), .O(n11836) );
  AOI22S U30100 ( .A1(n28913), .A2(n31532), .B1(n27919), .B2(img[1696]), .O(
        n28008) );
  ND2S U30101 ( .I1(n13819), .I2(img[1760]), .O(n28007) );
  ND3S U30102 ( .I1(n28425), .I2(n28008), .I3(n28007), .O(n28009) );
  AOI22S U30103 ( .A1(n28221), .A2(img[1760]), .B1(n13781), .B2(n31533), .O(
        n28010) );
  ND2S U30104 ( .I1(n28425), .I2(n28010), .O(n28011) );
  AOI22S U30105 ( .A1(n28075), .A2(n31534), .B1(n27919), .B2(img[1688]), .O(
        n28013) );
  AOI22S U30106 ( .A1(n13903), .A2(img[1752]), .B1(img[1784]), .B2(n13782), 
        .O(n28012) );
  ND3S U30107 ( .I1(n28425), .I2(n28013), .I3(n28012), .O(n28014) );
  MUX2 U30108 ( .A(img[1760]), .B(n28014), .S(n28933), .O(n11772) );
  AOI22S U30109 ( .A1(n28318), .A2(img[1784]), .B1(n13781), .B2(n31535), .O(
        n28015) );
  ND2S U30110 ( .I1(n28425), .I2(n28015), .O(n28016) );
  AOI22S U30111 ( .A1(n28075), .A2(n31536), .B1(n28069), .B2(img[1664]), .O(
        n28018) );
  AOI22S U30112 ( .A1(n13904), .A2(img[1728]), .B1(img[1760]), .B2(n28908), 
        .O(n28017) );
  ND3S U30113 ( .I1(n28425), .I2(n28018), .I3(n28017), .O(n28019) );
  MUX2 U30114 ( .A(img[1784]), .B(n28019), .S(n28941), .O(n11748) );
  AOI22S U30115 ( .A1(n26970), .A2(img[1728]), .B1(n28862), .B2(n31537), .O(
        n28020) );
  ND2S U30116 ( .I1(n28425), .I2(n28020), .O(n28021) );
  MUX2 U30117 ( .A(img[1720]), .B(n28021), .S(n28948), .O(n11812) );
  AOI22S U30118 ( .A1(n27735), .A2(n31538), .B1(n24313), .B2(img[1720]), .O(
        n28023) );
  ND3S U30119 ( .I1(n28425), .I2(n28023), .I3(n28022), .O(n28024) );
  MUX2 U30120 ( .A(img[1728]), .B(n28024), .S(n28945), .O(n11804) );
  AOI22S U30121 ( .A1(n13778), .A2(img[1624]), .B1(n13781), .B2(n31539), .O(
        n28025) );
  ND2S U30122 ( .I1(n28425), .I2(n28025), .O(n28026) );
  MUX2 U30123 ( .A(n28026), .B(img[1568]), .S(n28951), .O(n11964) );
  AOI22S U30124 ( .A1(n28075), .A2(n31540), .B1(n28069), .B2(img[1568]), .O(
        n28028) );
  ND2S U30125 ( .I1(n13820), .I2(img[1632]), .O(n28027) );
  ND3S U30126 ( .I1(n28425), .I2(n28028), .I3(n28027), .O(n28029) );
  AOI22S U30127 ( .A1(n28106), .A2(img[1632]), .B1(n13781), .B2(n31541), .O(
        n28030) );
  ND2S U30128 ( .I1(n28292), .I2(n28030), .O(n28031) );
  MUX2 U30129 ( .A(img[1560]), .B(n28031), .S(n28958), .O(n11972) );
  AOI22S U30130 ( .A1(n28075), .A2(n31542), .B1(n24313), .B2(img[1560]), .O(
        n28033) );
  AOI22S U30131 ( .A1(n13904), .A2(img[1624]), .B1(img[1656]), .B2(n13782), 
        .O(n28032) );
  ND3S U30132 ( .I1(n28425), .I2(n28033), .I3(n28032), .O(n28034) );
  MUX2 U30133 ( .A(img[1632]), .B(n28034), .S(n28962), .O(n11900) );
  AOI22S U30134 ( .A1(n28106), .A2(img[1656]), .B1(n28037), .B2(n31543), .O(
        n28035) );
  ND2S U30135 ( .I1(n28425), .I2(n28035), .O(n28036) );
  AOI22S U30136 ( .A1(n28037), .A2(n31544), .B1(n24313), .B2(img[1536]), .O(
        n28039) );
  AOI22S U30137 ( .A1(n13905), .A2(img[1600]), .B1(img[1632]), .B2(n13782), 
        .O(n28038) );
  ND3S U30138 ( .I1(n28425), .I2(n28039), .I3(n28038), .O(n28040) );
  MUX2 U30139 ( .A(img[1656]), .B(n28040), .S(n28969), .O(n11876) );
  AOI22S U30140 ( .A1(n28106), .A2(img[1600]), .B1(n27511), .B2(n31545), .O(
        n28041) );
  ND2S U30141 ( .I1(n28292), .I2(n28041), .O(n28042) );
  AOI22S U30142 ( .A1(n28075), .A2(n31546), .B1(n28069), .B2(img[1592]), .O(
        n28045) );
  ND3S U30143 ( .I1(n28425), .I2(n28045), .I3(n28044), .O(n28046) );
  MUX2 U30144 ( .A(img[1600]), .B(n28046), .S(n28973), .O(n11932) );
  AOI22S U30145 ( .A1(n28106), .A2(img[1144]), .B1(n25591), .B2(n31547), .O(
        n28047) );
  ND2S U30146 ( .I1(n28425), .I2(n28047), .O(n28048) );
  MUX2 U30147 ( .A(img[1024]), .B(n28048), .S(n28979), .O(n12508) );
  AOI22S U30148 ( .A1(n28162), .A2(n31548), .B1(n28069), .B2(img[1024]), .O(
        n28050) );
  ND2S U30149 ( .I1(n13820), .I2(img[1088]), .O(n28049) );
  ND3S U30150 ( .I1(n28425), .I2(n28050), .I3(n28049), .O(n28051) );
  MUX2 U30151 ( .A(img[1144]), .B(n28051), .S(n28983), .O(n12388) );
  AOI22S U30152 ( .A1(n13778), .A2(img[1088]), .B1(n13781), .B2(n31549), .O(
        n28052) );
  ND2S U30153 ( .I1(n28425), .I2(n28052), .O(n28053) );
  AOI22S U30154 ( .A1(n29397), .A2(n31550), .B1(n28069), .B2(img[1080]), .O(
        n28055) );
  ND2S U30155 ( .I1(n29124), .I2(img[1144]), .O(n28054) );
  ND3S U30156 ( .I1(n28425), .I2(n28055), .I3(n28054), .O(n28056) );
  MUX2 U30157 ( .A(img[1088]), .B(n28056), .S(n28987), .O(n12444) );
  AOI22S U30158 ( .A1(n13778), .A2(img[2008]), .B1(n29397), .B2(n31551), .O(
        n28057) );
  ND2S U30159 ( .I1(n28425), .I2(n28057), .O(n28058) );
  MUX2 U30160 ( .A(n28058), .B(img[1952]), .S(n28993), .O(n11580) );
  AOI22S U30161 ( .A1(n29242), .A2(n31552), .B1(n28069), .B2(img[1952]), .O(
        n28060) );
  ND3S U30162 ( .I1(n28425), .I2(n28060), .I3(n28059), .O(n28061) );
  AOI22S U30163 ( .A1(n13778), .A2(img[2016]), .B1(n25062), .B2(n31553), .O(
        n28062) );
  ND2S U30164 ( .I1(n28425), .I2(n28062), .O(n28063) );
  MUX2 U30165 ( .A(img[1944]), .B(n28063), .S(n29000), .O(n11588) );
  AOI22S U30166 ( .A1(n28182), .A2(n31554), .B1(n28069), .B2(img[1944]), .O(
        n28065) );
  AOI22S U30167 ( .A1(n13899), .A2(img[2008]), .B1(img[2040]), .B2(n13782), 
        .O(n28064) );
  ND3S U30168 ( .I1(n28425), .I2(n28065), .I3(n28064), .O(n28066) );
  MUX2 U30169 ( .A(img[2016]), .B(n28066), .S(n29004), .O(n11516) );
  AOI22S U30170 ( .A1(n13778), .A2(img[2040]), .B1(n13779), .B2(n31555), .O(
        n28067) );
  ND2S U30171 ( .I1(n28425), .I2(n28067), .O(n28068) );
  MUX2 U30172 ( .A(img[1920]), .B(n28068), .S(n29007), .O(n11612) );
  AOI22S U30173 ( .A1(n28075), .A2(n31556), .B1(n28069), .B2(img[1920]), .O(
        n28071) );
  AOI22S U30174 ( .A1(n13904), .A2(img[1984]), .B1(img[2016]), .B2(n13782), 
        .O(n28070) );
  ND3S U30175 ( .I1(n28425), .I2(n28071), .I3(n28070), .O(n28072) );
  AOI22S U30176 ( .A1(n13778), .A2(img[1984]), .B1(n28343), .B2(n31557), .O(
        n28073) );
  ND2S U30177 ( .I1(n28425), .I2(n28073), .O(n28074) );
  MUX2 U30178 ( .A(img[1976]), .B(n28074), .S(n29018), .O(n11556) );
  AOI22S U30179 ( .A1(n28075), .A2(n31558), .B1(n28254), .B2(img[1976]), .O(
        n28077) );
  ND2S U30180 ( .I1(n13820), .I2(img[2040]), .O(n28076) );
  ND3S U30181 ( .I1(n28425), .I2(n28077), .I3(n28076), .O(n28078) );
  MUX2 U30182 ( .A(img[1984]), .B(n28078), .S(n29015), .O(n11548) );
  AOI22S U30183 ( .A1(n13778), .A2(img[512]), .B1(n13781), .B2(n31559), .O(
        n28079) );
  ND2S U30184 ( .I1(n28292), .I2(n28079), .O(n28080) );
  AOI22S U30185 ( .A1(n13778), .A2(img[632]), .B1(n27049), .B2(n31560), .O(
        n28081) );
  ND2S U30186 ( .I1(n28425), .I2(n28081), .O(n28082) );
  AOI22S U30187 ( .A1(n28382), .A2(img[0]), .B1(n28614), .B2(n31561), .O(
        n28084) );
  ND2S U30188 ( .I1(n28425), .I2(n28084), .O(n28085) );
  MUX2 U30189 ( .A(img[120]), .B(n28085), .S(n29392), .O(n13412) );
  AOI22S U30190 ( .A1(n28382), .A2(img[120]), .B1(n25377), .B2(n31562), .O(
        n28086) );
  ND2S U30191 ( .I1(n28425), .I2(n28086), .O(n28087) );
  AOI22S U30192 ( .A1(n13773), .A2(img[896]), .B1(n28862), .B2(n31563), .O(
        n28088) );
  ND2S U30193 ( .I1(n28292), .I2(n28088), .O(n28089) );
  AOI22S U30194 ( .A1(n26822), .A2(img[1016]), .B1(n28614), .B2(n31564), .O(
        n28090) );
  ND2S U30195 ( .I1(n28425), .I2(n28090), .O(n28091) );
  AOI22S U30196 ( .A1(n28106), .A2(img[128]), .B1(n27049), .B2(n31565), .O(
        n28092) );
  ND2S U30197 ( .I1(n28425), .I2(n28092), .O(n28093) );
  MUX2 U30198 ( .A(img[248]), .B(n28093), .S(n29405), .O(n13284) );
  AOI22S U30199 ( .A1(n28106), .A2(img[248]), .B1(n28614), .B2(n31566), .O(
        n28094) );
  ND2S U30200 ( .I1(n28425), .I2(n28094), .O(n28095) );
  MUX2 U30201 ( .A(n28095), .B(img[128]), .S(n29402), .O(n13404) );
  AOI22S U30202 ( .A1(n28106), .A2(img[256]), .B1(n28614), .B2(n31567), .O(
        n28096) );
  ND2S U30203 ( .I1(n28425), .I2(n28096), .O(n28097) );
  MUX2 U30204 ( .A(img[376]), .B(n28097), .S(n29412), .O(n13156) );
  AOI22S U30205 ( .A1(n28106), .A2(img[376]), .B1(n28614), .B2(n31568), .O(
        n28098) );
  ND2S U30206 ( .I1(n28425), .I2(n28098), .O(n28099) );
  INV1S U30207 ( .I(img[504]), .O(n28100) );
  AOI22S U30208 ( .A1(n28106), .A2(img[384]), .B1(n28614), .B2(n28100), .O(
        n28101) );
  ND2S U30209 ( .I1(n28425), .I2(n28101), .O(n28102) );
  AOI22S U30210 ( .A1(n28106), .A2(img[504]), .B1(n29407), .B2(n31569), .O(
        n28103) );
  ND2S U30211 ( .I1(n28425), .I2(n28103), .O(n28104) );
  MUX2 U30212 ( .A(n28104), .B(img[384]), .S(n29416), .O(n13148) );
  INV1S U30213 ( .I(img[888]), .O(n28105) );
  AOI22S U30214 ( .A1(n28106), .A2(img[768]), .B1(n28614), .B2(n28105), .O(
        n28107) );
  ND2S U30215 ( .I1(n28425), .I2(n28107), .O(n28108) );
  AOI22S U30216 ( .A1(n27746), .A2(img[888]), .B1(n28614), .B2(n31570), .O(
        n28109) );
  ND2S U30217 ( .I1(n28425), .I2(n28109), .O(n28110) );
  MUX2 U30218 ( .A(img[768]), .B(n28110), .S(n29423), .O(n12764) );
  AOI22S U30219 ( .A1(n27746), .A2(img[640]), .B1(n28614), .B2(n31571), .O(
        n28111) );
  ND2S U30220 ( .I1(n28425), .I2(n28111), .O(n28112) );
  AOI22S U30221 ( .A1(n28083), .A2(img[760]), .B1(n28614), .B2(n31572), .O(
        n28113) );
  ND2S U30222 ( .I1(n28425), .I2(n28113), .O(n28114) );
  AOI22S U30223 ( .A1(n26822), .A2(img[616]), .B1(n29457), .B2(n31573), .O(
        n28115) );
  ND2S U30224 ( .I1(n13808), .I2(n28115), .O(n28116) );
  AOI22S U30225 ( .A1(n28083), .A2(img[528]), .B1(n28862), .B2(n31574), .O(
        n28117) );
  ND2S U30226 ( .I1(n13808), .I2(n28117), .O(n28118) );
  MUX2 U30227 ( .A(n28118), .B(img[616]), .S(n29024), .O(n12916) );
  AOI22S U30228 ( .A1(n29414), .A2(img[104]), .B1(n24193), .B2(n31575), .O(
        n28119) );
  ND2S U30229 ( .I1(n13808), .I2(n28119), .O(n28120) );
  MUX2 U30230 ( .A(img[16]), .B(n28120), .S(n29027), .O(n13516) );
  AOI22S U30231 ( .A1(n28083), .A2(img[16]), .B1(n23941), .B2(n31576), .O(
        n28121) );
  ND2S U30232 ( .I1(n13808), .I2(n28121), .O(n28122) );
  AOI22S U30233 ( .A1(n27990), .A2(img[1232]), .B1(n28862), .B2(n31577), .O(
        n28123) );
  ND2S U30234 ( .I1(n13808), .I2(n28123), .O(n28124) );
  MUX2 U30235 ( .A(img[1192]), .B(n28124), .S(n29033), .O(n12340) );
  AOI22S U30236 ( .A1(n28182), .A2(n31578), .B1(n28254), .B2(img[1192]), .O(
        n28126) );
  ND3S U30237 ( .I1(n28425), .I2(n28126), .I3(n28125), .O(n28127) );
  MUX2 U30238 ( .A(img[1232]), .B(n28127), .S(n29037), .O(n12300) );
  AOI22S U30239 ( .A1(n29414), .A2(img[1256]), .B1(n13781), .B2(n31579), .O(
        n28128) );
  ND2S U30240 ( .I1(n13808), .I2(n28128), .O(n28129) );
  AOI22S U30241 ( .A1(n25377), .A2(n31580), .B1(n28254), .B2(img[1168]), .O(
        n28131) );
  ND2S U30242 ( .I1(n29124), .I2(img[1232]), .O(n28130) );
  ND3S U30243 ( .I1(n28425), .I2(n28131), .I3(n28130), .O(n28132) );
  MUX2 U30244 ( .A(img[1256]), .B(n28132), .S(n29044), .O(n12276) );
  AOI22S U30245 ( .A1(n26822), .A2(img[1360]), .B1(n29407), .B2(n31581), .O(
        n28133) );
  ND2S U30246 ( .I1(n13808), .I2(n28133), .O(n28134) );
  MUX2 U30247 ( .A(n28134), .B(img[1320]), .S(n29047), .O(n12212) );
  AOI22S U30248 ( .A1(n28135), .A2(n31582), .B1(n28254), .B2(img[1320]), .O(
        n28137) );
  ND3S U30249 ( .I1(n28425), .I2(n28137), .I3(n28136), .O(n28138) );
  MUX2 U30250 ( .A(img[1360]), .B(n28138), .S(n29051), .O(n12172) );
  AOI22S U30251 ( .A1(n13773), .A2(img[1384]), .B1(n29194), .B2(n31583), .O(
        n28139) );
  ND2S U30252 ( .I1(n13808), .I2(n28139), .O(n28140) );
  MUX2 U30253 ( .A(n28140), .B(img[1296]), .S(n29054), .O(n12236) );
  AOI22S U30254 ( .A1(n28182), .A2(n31584), .B1(n28254), .B2(img[1296]), .O(
        n28142) );
  ND2S U30255 ( .I1(n13770), .I2(img[1360]), .O(n28141) );
  ND3S U30256 ( .I1(n28425), .I2(n28142), .I3(n28141), .O(n28143) );
  MUX2 U30257 ( .A(img[1384]), .B(n28143), .S(n29058), .O(n12148) );
  AOI22S U30258 ( .A1(n29414), .A2(img[1000]), .B1(n28862), .B2(n31585), .O(
        n28144) );
  ND2S U30259 ( .I1(n13808), .I2(n28144), .O(n28145) );
  MUX2 U30260 ( .A(img[912]), .B(n28145), .S(n29061), .O(n12620) );
  AOI22S U30261 ( .A1(n27987), .A2(img[912]), .B1(n13775), .B2(n31586), .O(
        n28146) );
  ND2S U30262 ( .I1(n13808), .I2(n28146), .O(n28147) );
  AOI22S U30263 ( .A1(n13776), .A2(img[232]), .B1(n28862), .B2(n31587), .O(
        n28148) );
  ND2S U30264 ( .I1(n13808), .I2(n28148), .O(n28149) );
  MUX2 U30265 ( .A(img[144]), .B(n28149), .S(n29067), .O(n13388) );
  AOI22S U30266 ( .A1(n25595), .A2(img[144]), .B1(n13781), .B2(n31588), .O(
        n28150) );
  ND2S U30267 ( .I1(n13808), .I2(n28150), .O(n28151) );
  MUX2 U30268 ( .A(img[232]), .B(n28151), .S(n29070), .O(n13300) );
  AOI22S U30269 ( .A1(n29414), .A2(img[360]), .B1(n13779), .B2(n31589), .O(
        n28152) );
  ND2S U30270 ( .I1(n13808), .I2(n28152), .O(n28153) );
  AOI22S U30271 ( .A1(n28382), .A2(img[272]), .B1(n24374), .B2(n31590), .O(
        n28154) );
  ND2S U30272 ( .I1(n13808), .I2(n28154), .O(n28155) );
  MUX2 U30273 ( .A(img[360]), .B(n28155), .S(n29078), .O(n13172) );
  AOI22S U30274 ( .A1(n27746), .A2(img[488]), .B1(n24374), .B2(n31591), .O(
        n28156) );
  ND2S U30275 ( .I1(n13808), .I2(n28156), .O(n28157) );
  AOI22S U30276 ( .A1(n28083), .A2(img[400]), .B1(n24374), .B2(n31592), .O(
        n28158) );
  ND2S U30277 ( .I1(n13808), .I2(n28158), .O(n28159) );
  MUX2 U30278 ( .A(img[488]), .B(n28159), .S(n29084), .O(n13044) );
  AOI22S U30279 ( .A1(n28347), .A2(img[1488]), .B1(n24374), .B2(n31593), .O(
        n28160) );
  ND2S U30280 ( .I1(n13808), .I2(n28160), .O(n28161) );
  MUX2 U30281 ( .A(n28161), .B(img[1448]), .S(n29087), .O(n12084) );
  AOI22S U30282 ( .A1(n28162), .A2(n31594), .B1(n24313), .B2(img[1448]), .O(
        n28164) );
  ND2S U30283 ( .I1(n13900), .I2(img[1512]), .O(n28163) );
  ND3S U30284 ( .I1(n28425), .I2(n28164), .I3(n28163), .O(n28165) );
  MUX2 U30285 ( .A(n28165), .B(img[1488]), .S(n29091), .O(n12044) );
  AOI22S U30286 ( .A1(n29414), .A2(img[1512]), .B1(n24374), .B2(n31595), .O(
        n28166) );
  ND2S U30287 ( .I1(n13808), .I2(n28166), .O(n28167) );
  MUX2 U30288 ( .A(img[1424]), .B(n28167), .S(n29094), .O(n12108) );
  AOI22S U30289 ( .A1(n28182), .A2(n31596), .B1(n28043), .B2(img[1424]), .O(
        n28169) );
  ND3S U30290 ( .I1(n28425), .I2(n28169), .I3(n28168), .O(n28170) );
  AOI22S U30291 ( .A1(n13773), .A2(img[872]), .B1(n24374), .B2(n31597), .O(
        n28171) );
  ND2S U30292 ( .I1(n13808), .I2(n28171), .O(n28172) );
  MUX2 U30293 ( .A(img[784]), .B(n28172), .S(n29102), .O(n12748) );
  INV1S U30294 ( .I(img[872]), .O(n28173) );
  AOI22S U30295 ( .A1(n13777), .A2(img[784]), .B1(n24374), .B2(n28173), .O(
        n28174) );
  ND2S U30296 ( .I1(n13808), .I2(n28174), .O(n28175) );
  AOI22S U30297 ( .A1(n13777), .A2(img[744]), .B1(n24374), .B2(n31598), .O(
        n28176) );
  ND2S U30298 ( .I1(n13808), .I2(n28176), .O(n28177) );
  AOI22S U30299 ( .A1(n13772), .A2(img[656]), .B1(n29530), .B2(n31599), .O(
        n28178) );
  ND2S U30300 ( .I1(n13808), .I2(n28178), .O(n28179) );
  MUX2 U30301 ( .A(n28179), .B(img[744]), .S(n29112), .O(n12788) );
  AOI22S U30302 ( .A1(n13780), .A2(img[1864]), .B1(n28433), .B2(n31600), .O(
        n28180) );
  ND2S U30303 ( .I1(n13808), .I2(n28180), .O(n28181) );
  MUX2 U30304 ( .A(n28181), .B(img[1840]), .S(n28693), .O(n11692) );
  AOI22S U30305 ( .A1(n28182), .A2(n31601), .B1(n24313), .B2(img[1840]), .O(
        n28184) );
  ND3S U30306 ( .I1(n28425), .I2(n28184), .I3(n28183), .O(n28185) );
  MUX2 U30307 ( .A(img[1864]), .B(n28185), .S(n28698), .O(n11668) );
  AOI22S U30308 ( .A1(n27990), .A2(img[1904]), .B1(n28614), .B2(n31602), .O(
        n28186) );
  ND2S U30309 ( .I1(n13808), .I2(n28186), .O(n28187) );
  AOI22S U30310 ( .A1(n25591), .A2(n31603), .B1(n28069), .B2(img[1800]), .O(
        n28189) );
  AOI22S U30311 ( .A1(n13899), .A2(img[1864]), .B1(img[1896]), .B2(n13782), 
        .O(n28188) );
  ND3S U30312 ( .I1(n28425), .I2(n28189), .I3(n28188), .O(n28190) );
  MUX2 U30313 ( .A(img[1904]), .B(n28190), .S(n28690), .O(n11628) );
  AOI22S U30314 ( .A1(n27065), .A2(img[1872]), .B1(n29397), .B2(n31604), .O(
        n28191) );
  ND2S U30315 ( .I1(n13808), .I2(n28191), .O(n28192) );
  MUX2 U30316 ( .A(n28192), .B(img[1832]), .S(n28672), .O(n11700) );
  AOI22S U30317 ( .A1(n28037), .A2(n31605), .B1(n24313), .B2(img[1832]), .O(
        n28194) );
  ND2S U30318 ( .I1(n13819), .I2(img[1896]), .O(n28193) );
  ND3S U30319 ( .I1(n28425), .I2(n28194), .I3(n28193), .O(n28195) );
  MUX2 U30320 ( .A(img[1872]), .B(n28195), .S(n28676), .O(n11660) );
  AOI22S U30321 ( .A1(n25810), .A2(img[1896]), .B1(n28135), .B2(n31606), .O(
        n28196) );
  ND2S U30322 ( .I1(n13808), .I2(n28196), .O(n28197) );
  AOI22S U30323 ( .A1(n28938), .A2(n31607), .B1(n28069), .B2(img[1808]), .O(
        n28199) );
  AOI22S U30324 ( .A1(n13905), .A2(img[1872]), .B1(img[1904]), .B2(n13782), 
        .O(n28198) );
  ND3S U30325 ( .I1(n28425), .I2(n28199), .I3(n28198), .O(n28200) );
  MUX2 U30326 ( .A(img[1896]), .B(n28200), .S(n28683), .O(n11636) );
  AOI22S U30327 ( .A1(n29072), .A2(img[1736]), .B1(n28614), .B2(n31608), .O(
        n28201) );
  ND2S U30328 ( .I1(n28292), .I2(n28201), .O(n28202) );
  AOI22S U30329 ( .A1(n28695), .A2(n31609), .B1(n28069), .B2(img[1712]), .O(
        n28204) );
  ND2S U30330 ( .I1(n13905), .I2(img[1776]), .O(n28203) );
  AOI22S U30331 ( .A1(n26490), .A2(img[1776]), .B1(n29096), .B2(n31610), .O(
        n28206) );
  ND2S U30332 ( .I1(n28292), .I2(n28206), .O(n28207) );
  MUX2 U30333 ( .A(img[1672]), .B(n28207), .S(n28715), .O(n11860) );
  AOI22S U30334 ( .A1(n28075), .A2(n31611), .B1(n28069), .B2(img[1672]), .O(
        n28209) );
  AOI22S U30335 ( .A1(n13820), .A2(img[1736]), .B1(img[1768]), .B2(n13782), 
        .O(n28208) );
  ND3S U30336 ( .I1(n28425), .I2(n28209), .I3(n28208), .O(n28210) );
  MUX2 U30337 ( .A(img[1776]), .B(n28210), .S(n28719), .O(n11756) );
  AOI22S U30338 ( .A1(n27685), .A2(img[1744]), .B1(n29407), .B2(n31612), .O(
        n28211) );
  ND2S U30339 ( .I1(n28292), .I2(n28211), .O(n28212) );
  AOI22S U30340 ( .A1(n28182), .A2(n31613), .B1(n28069), .B2(img[1704]), .O(
        n28214) );
  ND2S U30341 ( .I1(n13770), .I2(img[1768]), .O(n28213) );
  ND3S U30342 ( .I1(n28425), .I2(n28214), .I3(n28213), .O(n28215) );
  MUX2 U30343 ( .A(img[1744]), .B(n28215), .S(n28705), .O(n11788) );
  AOI22S U30344 ( .A1(n25810), .A2(img[1768]), .B1(n28433), .B2(n31614), .O(
        n28216) );
  ND2S U30345 ( .I1(n28292), .I2(n28216), .O(n28217) );
  AOI22S U30346 ( .A1(n25377), .A2(n31615), .B1(n28254), .B2(img[1680]), .O(
        n28219) );
  AOI22S U30347 ( .A1(n13905), .A2(img[1744]), .B1(img[1776]), .B2(n13782), 
        .O(n28218) );
  ND3S U30348 ( .I1(n28425), .I2(n28219), .I3(n28218), .O(n28220) );
  MUX2 U30349 ( .A(img[1768]), .B(n28220), .S(n28712), .O(n11764) );
  AOI22S U30350 ( .A1(n29129), .A2(img[1608]), .B1(n29096), .B2(n31616), .O(
        n28222) );
  ND2S U30351 ( .I1(n28292), .I2(n28222), .O(n28223) );
  AOI22S U30352 ( .A1(n28135), .A2(n31617), .B1(n28254), .B2(img[1584]), .O(
        n28225) );
  ND3S U30353 ( .I1(n28425), .I2(n28225), .I3(n28224), .O(n28226) );
  MUX2 U30354 ( .A(img[1608]), .B(n28226), .S(n28754), .O(n11924) );
  AOI22S U30355 ( .A1(n28106), .A2(img[1648]), .B1(n29530), .B2(n31618), .O(
        n28227) );
  ND2S U30356 ( .I1(n28292), .I2(n28227), .O(n28228) );
  AOI22S U30357 ( .A1(n28614), .A2(n31619), .B1(n28254), .B2(img[1544]), .O(
        n28230) );
  AOI22S U30358 ( .A1(n29124), .A2(img[1608]), .B1(img[1640]), .B2(n13782), 
        .O(n28229) );
  ND3S U30359 ( .I1(n28425), .I2(n28230), .I3(n28229), .O(n28231) );
  MUX2 U30360 ( .A(img[1648]), .B(n28231), .S(n28747), .O(n11884) );
  AOI22S U30361 ( .A1(n25595), .A2(img[1616]), .B1(n29530), .B2(n31620), .O(
        n28232) );
  ND2S U30362 ( .I1(n28292), .I2(n28232), .O(n28233) );
  AOI22S U30363 ( .A1(n28938), .A2(n31621), .B1(n28254), .B2(img[1576]), .O(
        n28235) );
  ND3S U30364 ( .I1(n28425), .I2(n28235), .I3(n28234), .O(n28236) );
  MUX2 U30365 ( .A(img[1616]), .B(n28236), .S(n28733), .O(n11916) );
  AOI22S U30366 ( .A1(n26855), .A2(img[1640]), .B1(n28614), .B2(n31622), .O(
        n28237) );
  ND2S U30367 ( .I1(n28292), .I2(n28237), .O(n28238) );
  AOI22S U30368 ( .A1(n28938), .A2(n31623), .B1(n28254), .B2(img[1552]), .O(
        n28240) );
  AOI22S U30369 ( .A1(n29124), .A2(img[1616]), .B1(img[1648]), .B2(n13782), 
        .O(n28239) );
  ND3S U30370 ( .I1(n28425), .I2(n28240), .I3(n28239), .O(n28241) );
  MUX2 U30371 ( .A(img[1640]), .B(n28241), .S(n28740), .O(n11892) );
  AOI22S U30372 ( .A1(n28840), .A2(img[1104]), .B1(n24374), .B2(n31624), .O(
        n28242) );
  ND2S U30373 ( .I1(n28292), .I2(n28242), .O(n28243) );
  AOI22S U30374 ( .A1(n28182), .A2(n31625), .B1(n28254), .B2(img[1064]), .O(
        n28245) );
  ND2S U30375 ( .I1(n29124), .I2(img[1128]), .O(n28244) );
  ND3S U30376 ( .I1(n28425), .I2(n28245), .I3(n28244), .O(n28246) );
  MUX2 U30377 ( .A(img[1104]), .B(n28246), .S(n29119), .O(n12428) );
  AOI22S U30378 ( .A1(n13771), .A2(img[1128]), .B1(n13779), .B2(n31626), .O(
        n28247) );
  ND2S U30379 ( .I1(n28292), .I2(n28247), .O(n28248) );
  AOI22S U30380 ( .A1(n28938), .A2(n31627), .B1(n28254), .B2(img[1040]), .O(
        n28250) );
  ND2S U30381 ( .I1(n29124), .I2(img[1104]), .O(n28249) );
  ND3S U30382 ( .I1(n28425), .I2(n28250), .I3(n28249), .O(n28251) );
  MUX2 U30383 ( .A(img[1128]), .B(n28251), .S(n29127), .O(n12404) );
  AOI22S U30384 ( .A1(n13772), .A2(img[1992]), .B1(n28343), .B2(n31628), .O(
        n28252) );
  ND2S U30385 ( .I1(n28292), .I2(n28252), .O(n28253) );
  AOI22S U30386 ( .A1(n28135), .A2(n31629), .B1(n28254), .B2(img[1968]), .O(
        n28256) );
  ND2S U30387 ( .I1(n29124), .I2(img[2032]), .O(n28255) );
  ND3S U30388 ( .I1(n28425), .I2(n28256), .I3(n28255), .O(n28257) );
  MUX2 U30389 ( .A(img[1992]), .B(n28257), .S(n28796), .O(n11540) );
  AOI22S U30390 ( .A1(n13771), .A2(img[2032]), .B1(n29194), .B2(n31630), .O(
        n28258) );
  ND2S U30391 ( .I1(n28292), .I2(n28258), .O(n28259) );
  MUX2 U30392 ( .A(img[1928]), .B(n28259), .S(n28785), .O(n11604) );
  AOI22S U30393 ( .A1(n24193), .A2(n31631), .B1(n28069), .B2(img[1928]), .O(
        n28261) );
  AOI22S U30394 ( .A1(n29124), .A2(img[1992]), .B1(img[2024]), .B2(n13782), 
        .O(n28260) );
  ND3S U30395 ( .I1(n28425), .I2(n28261), .I3(n28260), .O(n28262) );
  MUX2 U30396 ( .A(img[2032]), .B(n28262), .S(n28789), .O(n11500) );
  AOI22S U30397 ( .A1(n13778), .A2(img[2000]), .B1(n24374), .B2(n31632), .O(
        n28263) );
  ND2S U30398 ( .I1(n28292), .I2(n28263), .O(n28264) );
  AOI22S U30399 ( .A1(n28938), .A2(n31633), .B1(n24313), .B2(img[1960]), .O(
        n28266) );
  ND2S U30400 ( .I1(n13903), .I2(img[2024]), .O(n28265) );
  ND3S U30401 ( .I1(n28425), .I2(n28266), .I3(n28265), .O(n28267) );
  MUX2 U30402 ( .A(img[2000]), .B(n28267), .S(n28775), .O(n11532) );
  AOI22S U30403 ( .A1(n13777), .A2(img[2024]), .B1(n13781), .B2(n31634), .O(
        n28268) );
  ND2S U30404 ( .I1(n28292), .I2(n28268), .O(n28269) );
  AOI22S U30405 ( .A1(n28938), .A2(n31635), .B1(n28043), .B2(img[1936]), .O(
        n28271) );
  AOI22S U30406 ( .A1(n13904), .A2(img[2000]), .B1(img[2032]), .B2(n13782), 
        .O(n28270) );
  ND3S U30407 ( .I1(n28425), .I2(n28271), .I3(n28270), .O(n28272) );
  MUX2 U30408 ( .A(img[2024]), .B(n28272), .S(n28782), .O(n11508) );
  AOI22S U30409 ( .A1(n13780), .A2(img[520]), .B1(n25591), .B2(n31636), .O(
        n28273) );
  ND2S U30410 ( .I1(n28292), .I2(n28273), .O(n28274) );
  AOI22S U30411 ( .A1(n28318), .A2(img[624]), .B1(n25062), .B2(n31637), .O(
        n28275) );
  ND2S U30412 ( .I1(n28292), .I2(n28275), .O(n28276) );
  AOI22S U30413 ( .A1(n13776), .A2(img[8]), .B1(n28433), .B2(n31638), .O(
        n28277) );
  ND2S U30414 ( .I1(n28292), .I2(n28277), .O(n28278) );
  MUX2 U30415 ( .A(img[112]), .B(n28278), .S(n29536), .O(n13420) );
  AOI22S U30416 ( .A1(n29076), .A2(img[112]), .B1(n28862), .B2(n31639), .O(
        n28279) );
  ND2S U30417 ( .I1(n28292), .I2(n28279), .O(n28280) );
  AOI22S U30418 ( .A1(n29129), .A2(img[1224]), .B1(n28343), .B2(n31640), .O(
        n28281) );
  ND2S U30419 ( .I1(n28292), .I2(n28281), .O(n28282) );
  AOI22S U30420 ( .A1(n28938), .A2(n31641), .B1(n28043), .B2(img[1200]), .O(
        n28284) );
  ND3S U30421 ( .I1(n28425), .I2(n28284), .I3(n28283), .O(n28285) );
  MUX2 U30422 ( .A(img[1224]), .B(n28285), .S(n28602), .O(n12308) );
  AOI22S U30423 ( .A1(n28938), .A2(n31642), .B1(n24946), .B2(img[1160]), .O(
        n28287) );
  ND3S U30424 ( .I1(n28425), .I2(n28287), .I3(n28286), .O(n28288) );
  MUX2 U30425 ( .A(img[1264]), .B(n28288), .S(n28595), .O(n12268) );
  AOI22S U30426 ( .A1(n28347), .A2(img[1264]), .B1(n28343), .B2(n31643), .O(
        n28289) );
  ND2S U30427 ( .I1(n28292), .I2(n28289), .O(n28290) );
  AOI22S U30428 ( .A1(n13772), .A2(img[1352]), .B1(n23918), .B2(n31644), .O(
        n28291) );
  ND2S U30429 ( .I1(n28292), .I2(n28291), .O(n28293) );
  AOI22S U30430 ( .A1(n28614), .A2(n31645), .B1(n24313), .B2(img[1328]), .O(
        n28295) );
  ND3S U30431 ( .I1(n28425), .I2(n28295), .I3(n28294), .O(n28296) );
  MUX2 U30432 ( .A(img[1352]), .B(n28296), .S(n28617), .O(n12180) );
  AOI22S U30433 ( .A1(n25062), .A2(n31646), .B1(n24313), .B2(img[1288]), .O(
        n28298) );
  ND2S U30434 ( .I1(n13770), .I2(img[1352]), .O(n28297) );
  ND3S U30435 ( .I1(n28425), .I2(n28298), .I3(n28297), .O(n28299) );
  MUX2 U30436 ( .A(img[1392]), .B(n28299), .S(n28609), .O(n12140) );
  AOI22S U30437 ( .A1(n28347), .A2(img[1392]), .B1(n25062), .B2(n31647), .O(
        n28300) );
  ND2S U30438 ( .I1(n28425), .I2(n28300), .O(n28301) );
  AOI22S U30439 ( .A1(n28221), .A2(img[904]), .B1(n28135), .B2(n31648), .O(
        n28302) );
  ND2S U30440 ( .I1(n28425), .I2(n28302), .O(n28303) );
  MUX2 U30441 ( .A(img[1008]), .B(n28303), .S(n29303), .O(n12524) );
  AOI22S U30442 ( .A1(n29435), .A2(img[1008]), .B1(n28433), .B2(n31649), .O(
        n28304) );
  ND2S U30443 ( .I1(n28425), .I2(n28304), .O(n28305) );
  AOI22S U30444 ( .A1(n28840), .A2(img[136]), .B1(n28343), .B2(n31650), .O(
        n28306) );
  ND2S U30445 ( .I1(n28425), .I2(n28306), .O(n28307) );
  MUX2 U30446 ( .A(img[240]), .B(n28307), .S(n29309), .O(n13292) );
  AOI22S U30447 ( .A1(n13771), .A2(img[240]), .B1(n28862), .B2(n31651), .O(
        n28308) );
  ND2S U30448 ( .I1(n28425), .I2(n28308), .O(n28309) );
  AOI22S U30449 ( .A1(n29076), .A2(img[264]), .B1(n29530), .B2(n31652), .O(
        n28310) );
  ND2S U30450 ( .I1(n28425), .I2(n28310), .O(n28311) );
  AOI22S U30451 ( .A1(n29076), .A2(img[368]), .B1(n25591), .B2(n31653), .O(
        n28312) );
  ND2S U30452 ( .I1(n28425), .I2(n28312), .O(n28313) );
  MUX2 U30453 ( .A(n28313), .B(img[264]), .S(n29312), .O(n13268) );
  AOI22S U30454 ( .A1(n29076), .A2(img[392]), .B1(n29407), .B2(n31654), .O(
        n28314) );
  ND2S U30455 ( .I1(n28425), .I2(n28314), .O(n28315) );
  AOI22S U30456 ( .A1(n26970), .A2(img[496]), .B1(n13775), .B2(n31655), .O(
        n28316) );
  ND2S U30457 ( .I1(n28425), .I2(n28316), .O(n28317) );
  AOI22S U30458 ( .A1(n29414), .A2(img[1480]), .B1(n28343), .B2(n31656), .O(
        n28319) );
  ND2S U30459 ( .I1(n28425), .I2(n28319), .O(n28320) );
  AOI22S U30460 ( .A1(n28938), .A2(n31657), .B1(n24313), .B2(img[1456]), .O(
        n28322) );
  ND3S U30461 ( .I1(n28425), .I2(n28322), .I3(n28321), .O(n28323) );
  MUX2 U30462 ( .A(img[1480]), .B(n28323), .S(n28656), .O(n12052) );
  AOI22S U30463 ( .A1(n28614), .A2(n31658), .B1(n24313), .B2(img[1416]), .O(
        n28325) );
  ND3S U30464 ( .I1(n28425), .I2(n28325), .I3(n28324), .O(n28326) );
  AOI22S U30465 ( .A1(n28347), .A2(img[1520]), .B1(n24193), .B2(n31659), .O(
        n28327) );
  ND2S U30466 ( .I1(n28292), .I2(n28327), .O(n28328) );
  INV1S U30467 ( .I(img[880]), .O(n28329) );
  AOI22S U30468 ( .A1(n28318), .A2(img[776]), .B1(n29407), .B2(n28329), .O(
        n28330) );
  ND2S U30469 ( .I1(n28425), .I2(n28330), .O(n28331) );
  AOI22S U30470 ( .A1(n28840), .A2(img[880]), .B1(n25591), .B2(n31660), .O(
        n28332) );
  ND2S U30471 ( .I1(n28425), .I2(n28332), .O(n28333) );
  MUX2 U30472 ( .A(img[776]), .B(n28333), .S(n29324), .O(n12756) );
  AOI22S U30473 ( .A1(n26822), .A2(img[648]), .B1(n25591), .B2(n31661), .O(
        n28334) );
  ND2S U30474 ( .I1(n28425), .I2(n28334), .O(n28335) );
  AOI22S U30475 ( .A1(n28347), .A2(img[752]), .B1(n29457), .B2(n31662), .O(
        n28336) );
  ND2S U30476 ( .I1(n28292), .I2(n28336), .O(n28337) );
  AOI22S U30477 ( .A1(n28382), .A2(img[1096]), .B1(n25591), .B2(n31663), .O(
        n28338) );
  ND2S U30478 ( .I1(n28425), .I2(n28338), .O(n28339) );
  AOI22S U30479 ( .A1(n25062), .A2(n31664), .B1(n28069), .B2(img[1072]), .O(
        n28341) );
  ND2S U30480 ( .I1(n13901), .I2(img[1136]), .O(n28340) );
  ND3S U30481 ( .I1(n28425), .I2(n28341), .I3(n28340), .O(n28342) );
  MUX2 U30482 ( .A(img[1096]), .B(n28342), .S(n28768), .O(n12436) );
  AOI22S U30483 ( .A1(n28343), .A2(n31665), .B1(n28043), .B2(img[1032]), .O(
        n28345) );
  ND2S U30484 ( .I1(n29124), .I2(img[1096]), .O(n28344) );
  ND3S U30485 ( .I1(n28425), .I2(n28345), .I3(n28344), .O(n28346) );
  MUX2 U30486 ( .A(img[1136]), .B(n28346), .S(n28761), .O(n12396) );
  AOI22S U30487 ( .A1(n28347), .A2(img[1136]), .B1(n29397), .B2(n31666), .O(
        n28348) );
  ND2S U30488 ( .I1(n28425), .I2(n28348), .O(n28349) );
  AOI22S U30489 ( .A1(n28347), .A2(img[600]), .B1(n29457), .B2(n31667), .O(
        n28350) );
  ND2S U30490 ( .I1(n28425), .I2(n28350), .O(n28351) );
  AOI22S U30491 ( .A1(n28347), .A2(img[544]), .B1(n29397), .B2(n31668), .O(
        n28352) );
  ND2S U30492 ( .I1(n28425), .I2(n28352), .O(n28353) );
  MUX2 U30493 ( .A(n28353), .B(img[600]), .S(n29478), .O(n12932) );
  AOI22S U30494 ( .A1(n28347), .A2(img[88]), .B1(n25062), .B2(n31669), .O(
        n28354) );
  ND2S U30495 ( .I1(n28425), .I2(n28354), .O(n28355) );
  AOI22S U30496 ( .A1(n29076), .A2(img[32]), .B1(n13779), .B2(n31670), .O(
        n28356) );
  ND2S U30497 ( .I1(n28292), .I2(n28356), .O(n28357) );
  MUX2 U30498 ( .A(img[88]), .B(n28357), .S(n29339), .O(n13444) );
  AOI22S U30499 ( .A1(n29076), .A2(img[1248]), .B1(n13779), .B2(n31671), .O(
        n28358) );
  ND2S U30500 ( .I1(n28425), .I2(n28358), .O(n28359) );
  MUX2 U30501 ( .A(img[1176]), .B(n28359), .S(n29214), .O(n12356) );
  AOI22S U30502 ( .A1(n25062), .A2(n31672), .B1(n25444), .B2(img[1176]), .O(
        n28361) );
  ND3S U30503 ( .I1(n28425), .I2(n28361), .I3(n28360), .O(n28362) );
  MUX2 U30504 ( .A(img[1248]), .B(n28362), .S(n29218), .O(n12284) );
  AOI22S U30505 ( .A1(n29076), .A2(img[1240]), .B1(n13781), .B2(n31673), .O(
        n28363) );
  ND2S U30506 ( .I1(n28425), .I2(n28363), .O(n28364) );
  MUX2 U30507 ( .A(n28364), .B(img[1184]), .S(n29207), .O(n12348) );
  AOI22S U30508 ( .A1(n29242), .A2(n31674), .B1(n25444), .B2(img[1184]), .O(
        n28366) );
  ND2S U30509 ( .I1(n29124), .I2(img[1248]), .O(n28365) );
  ND3S U30510 ( .I1(n28425), .I2(n28366), .I3(n28365), .O(n28367) );
  MUX2 U30511 ( .A(img[1240]), .B(n28367), .S(n29211), .O(n12292) );
  AOI22S U30512 ( .A1(n29076), .A2(img[1376]), .B1(n28695), .B2(n31675), .O(
        n28368) );
  ND2S U30513 ( .I1(n28425), .I2(n28368), .O(n28369) );
  MUX2 U30514 ( .A(img[1304]), .B(n28369), .S(n29240), .O(n12228) );
  AOI22S U30515 ( .A1(n25062), .A2(n31676), .B1(n25444), .B2(img[1304]), .O(
        n28371) );
  ND2S U30516 ( .I1(n13770), .I2(img[1368]), .O(n28370) );
  ND3S U30517 ( .I1(n28425), .I2(n28371), .I3(n28370), .O(n28372) );
  MUX2 U30518 ( .A(img[1376]), .B(n28372), .S(n29245), .O(n12156) );
  AOI22S U30519 ( .A1(n29076), .A2(img[1368]), .B1(n29397), .B2(n31677), .O(
        n28373) );
  ND2S U30520 ( .I1(n28425), .I2(n28373), .O(n28374) );
  MUX2 U30521 ( .A(n28374), .B(img[1312]), .S(n29233), .O(n12220) );
  AOI22S U30522 ( .A1(n25062), .A2(n31678), .B1(n25444), .B2(img[1312]), .O(
        n28376) );
  ND2S U30523 ( .I1(n29124), .I2(img[1376]), .O(n28375) );
  ND3S U30524 ( .I1(n28425), .I2(n28376), .I3(n28375), .O(n28377) );
  MUX2 U30525 ( .A(img[1368]), .B(n28377), .S(n29237), .O(n12164) );
  AOI22S U30526 ( .A1(n29076), .A2(img[984]), .B1(n24193), .B2(n31679), .O(
        n28378) );
  ND2S U30527 ( .I1(n28425), .I2(n28378), .O(n28379) );
  AOI22S U30528 ( .A1(n29076), .A2(img[928]), .B1(n28862), .B2(n31680), .O(
        n28380) );
  ND2S U30529 ( .I1(n28425), .I2(n28380), .O(n28381) );
  BUF1 U30530 ( .I(n28382), .O(n28442) );
  AOI22S U30531 ( .A1(n28442), .A2(img[216]), .B1(n13779), .B2(n31681), .O(
        n28383) );
  ND2S U30532 ( .I1(n28292), .I2(n28383), .O(n28384) );
  MUX2 U30533 ( .A(img[160]), .B(n28384), .S(n29355), .O(n13372) );
  AOI22S U30534 ( .A1(n28442), .A2(img[160]), .B1(n25591), .B2(n31682), .O(
        n28385) );
  ND2S U30535 ( .I1(n28425), .I2(n28385), .O(n28386) );
  MUX2 U30536 ( .A(img[216]), .B(n28386), .S(n29351), .O(n13316) );
  AOI22S U30537 ( .A1(n28442), .A2(img[344]), .B1(n13781), .B2(n31683), .O(
        n28387) );
  ND2S U30538 ( .I1(n28292), .I2(n28387), .O(n28388) );
  AOI22S U30539 ( .A1(n28442), .A2(img[288]), .B1(n25468), .B2(n31684), .O(
        n28389) );
  ND2S U30540 ( .I1(n28292), .I2(n28389), .O(n28390) );
  MUX2 U30541 ( .A(img[344]), .B(n28390), .S(n29358), .O(n13188) );
  AOI22S U30542 ( .A1(n28347), .A2(img[472]), .B1(n28135), .B2(n31685), .O(
        n28391) );
  ND2S U30543 ( .I1(n28425), .I2(n28391), .O(n28392) );
  MUX2 U30544 ( .A(img[416]), .B(n28392), .S(n29367), .O(n13116) );
  AOI22S U30545 ( .A1(n28347), .A2(img[416]), .B1(n28075), .B2(n31686), .O(
        n28393) );
  ND2S U30546 ( .I1(n28425), .I2(n28393), .O(n28394) );
  AOI22S U30547 ( .A1(n28347), .A2(img[1504]), .B1(n28695), .B2(n31687), .O(
        n28395) );
  ND2S U30548 ( .I1(n28425), .I2(n28395), .O(n28396) );
  MUX2 U30549 ( .A(n28396), .B(img[1432]), .S(n29255), .O(n12100) );
  AOI22S U30550 ( .A1(n25062), .A2(n31688), .B1(n25444), .B2(img[1432]), .O(
        n28398) );
  ND3S U30551 ( .I1(n28425), .I2(n28398), .I3(n28397), .O(n28399) );
  MUX2 U30552 ( .A(img[1504]), .B(n28399), .S(n29261), .O(n12028) );
  AOI22S U30553 ( .A1(n28347), .A2(img[1496]), .B1(n28433), .B2(n31689), .O(
        n28400) );
  ND2S U30554 ( .I1(n28425), .I2(n28400), .O(n28401) );
  MUX2 U30555 ( .A(n28401), .B(img[1440]), .S(n29248), .O(n12092) );
  AOI22S U30556 ( .A1(n28592), .A2(n31690), .B1(n28069), .B2(img[1440]), .O(
        n28403) );
  ND3S U30557 ( .I1(n28425), .I2(n28403), .I3(n28402), .O(n28404) );
  AOI22S U30558 ( .A1(n28347), .A2(img[856]), .B1(n28433), .B2(n31691), .O(
        n28405) );
  ND2S U30559 ( .I1(n28425), .I2(n28405), .O(n28406) );
  MUX2 U30560 ( .A(n28406), .B(img[800]), .S(n29374), .O(n12732) );
  INV1S U30561 ( .I(img[856]), .O(n28407) );
  AOI22S U30562 ( .A1(n28347), .A2(img[800]), .B1(n28433), .B2(n28407), .O(
        n28408) );
  ND2S U30563 ( .I1(n28425), .I2(n28408), .O(n28409) );
  AOI22S U30564 ( .A1(n28347), .A2(img[728]), .B1(n28433), .B2(n31692), .O(
        n28410) );
  ND2S U30565 ( .I1(n28425), .I2(n28410), .O(n28411) );
  AOI22S U30566 ( .A1(n28106), .A2(img[672]), .B1(n28433), .B2(n31693), .O(
        n28413) );
  ND2S U30567 ( .I1(n28425), .I2(n28413), .O(n28414) );
  AOI22S U30568 ( .A1(n28840), .A2(img[1120]), .B1(n28433), .B2(n31694), .O(
        n28416) );
  ND2S U30569 ( .I1(n13808), .I2(n28416), .O(n28417) );
  AOI22S U30570 ( .A1(n28433), .A2(n31695), .B1(n28069), .B2(img[1048]), .O(
        n28419) );
  ND2S U30571 ( .I1(n29258), .I2(img[1112]), .O(n28418) );
  ND3S U30572 ( .I1(n28425), .I2(n28419), .I3(n28418), .O(n28420) );
  MUX2 U30573 ( .A(img[1120]), .B(n28420), .S(n29198), .O(n12412) );
  AOI22S U30574 ( .A1(n28382), .A2(img[1112]), .B1(n28433), .B2(n31696), .O(
        n28421) );
  ND2S U30575 ( .I1(n13808), .I2(n28421), .O(n28422) );
  AOI22S U30576 ( .A1(n28592), .A2(n31697), .B1(n24313), .B2(img[1056]), .O(
        n28424) );
  ND2S U30577 ( .I1(n13900), .I2(img[1120]), .O(n28423) );
  ND3S U30578 ( .I1(n28425), .I2(n28424), .I3(n28423), .O(n28426) );
  MUX2 U30579 ( .A(img[1112]), .B(n28426), .S(n29189), .O(n12420) );
  AOI22S U30580 ( .A1(n26855), .A2(img[208]), .B1(n28433), .B2(n31698), .O(
        n28427) );
  ND2S U30581 ( .I1(n13808), .I2(n28427), .O(n28428) );
  MUX2 U30582 ( .A(img[168]), .B(n28428), .S(n29148), .O(n13364) );
  AOI22S U30583 ( .A1(n28442), .A2(img[168]), .B1(n28433), .B2(n31699), .O(
        n28429) );
  ND2S U30584 ( .I1(n13808), .I2(n28429), .O(n28430) );
  MUX2 U30585 ( .A(img[208]), .B(n28430), .S(n29151), .O(n13324) );
  AOI22S U30586 ( .A1(n28442), .A2(img[552]), .B1(n28433), .B2(n31700), .O(
        n28431) );
  ND2S U30587 ( .I1(n13808), .I2(n28431), .O(n28432) );
  MUX2 U30588 ( .A(n28432), .B(img[592]), .S(n29133), .O(n12940) );
  AOI22S U30589 ( .A1(n28442), .A2(img[80]), .B1(n28433), .B2(n31701), .O(
        n28434) );
  ND2S U30590 ( .I1(n13808), .I2(n28434), .O(n28435) );
  MUX2 U30591 ( .A(img[40]), .B(n28435), .S(n29136), .O(n13492) );
  AOI22S U30592 ( .A1(n28442), .A2(img[40]), .B1(n24193), .B2(n31702), .O(
        n28436) );
  ND2S U30593 ( .I1(n13808), .I2(n28436), .O(n28437) );
  AOI22S U30594 ( .A1(n28442), .A2(img[976]), .B1(n25591), .B2(n31703), .O(
        n28438) );
  ND2S U30595 ( .I1(n13808), .I2(n28438), .O(n28439) );
  AOI22S U30596 ( .A1(n28442), .A2(img[936]), .B1(n25062), .B2(n31704), .O(
        n28440) );
  ND2S U30597 ( .I1(n13808), .I2(n28440), .O(n28441) );
  MUX2 U30598 ( .A(img[976]), .B(n28441), .S(n29145), .O(n12556) );
  AOI22S U30599 ( .A1(n28442), .A2(img[336]), .B1(n28862), .B2(n31705), .O(
        n28443) );
  ND2S U30600 ( .I1(n13808), .I2(n28443), .O(n28444) );
  AOI22S U30601 ( .A1(n28347), .A2(img[296]), .B1(n25859), .B2(n31706), .O(
        n28445) );
  ND2S U30602 ( .I1(n13808), .I2(n28445), .O(n28446) );
  MUX2 U30603 ( .A(img[336]), .B(n28446), .S(n29157), .O(n13196) );
  AOI22S U30604 ( .A1(n13780), .A2(img[464]), .B1(n13781), .B2(n31707), .O(
        n28447) );
  ND2S U30605 ( .I1(n13808), .I2(n28447), .O(n28448) );
  AOI22S U30606 ( .A1(n27746), .A2(img[424]), .B1(n28614), .B2(n31708), .O(
        n28449) );
  ND2S U30607 ( .I1(n13808), .I2(n28449), .O(n28450) );
  MUX2 U30608 ( .A(img[464]), .B(n28450), .S(n29163), .O(n13068) );
  AOI22S U30609 ( .A1(n28347), .A2(img[848]), .B1(n29397), .B2(n31709), .O(
        n28451) );
  ND2S U30610 ( .I1(n13808), .I2(n28451), .O(n28452) );
  MUX2 U30611 ( .A(n28452), .B(img[808]), .S(n29166), .O(n12724) );
  INV1S U30612 ( .I(img[848]), .O(n28453) );
  AOI22S U30613 ( .A1(n29435), .A2(img[808]), .B1(n13781), .B2(n28453), .O(
        n28454) );
  ND2S U30614 ( .I1(n13808), .I2(n28454), .O(n28455) );
  AOI22S U30615 ( .A1(n29435), .A2(img[720]), .B1(n29397), .B2(n31710), .O(
        n28456) );
  ND2S U30616 ( .I1(n13808), .I2(n28456), .O(n28457) );
  MUX2 U30617 ( .A(n28457), .B(img[680]), .S(n29173), .O(n12852) );
  AOI22S U30618 ( .A1(n13773), .A2(img[680]), .B1(n28162), .B2(n31711), .O(
        n28458) );
  ND2S U30619 ( .I1(n13808), .I2(n28458), .O(n28459) );
  AOI22S U30620 ( .A1(n26970), .A2(img[584]), .B1(n28182), .B2(n31712), .O(
        n28460) );
  ND2S U30621 ( .I1(n13808), .I2(n28460), .O(n28461) );
  MUX2 U30622 ( .A(n28461), .B(img[560]), .S(n28578), .O(n12972) );
  AOI22S U30623 ( .A1(n28442), .A2(img[560]), .B1(n28162), .B2(n31713), .O(
        n28462) );
  ND2S U30624 ( .I1(n13808), .I2(n28462), .O(n28463) );
  MUX2 U30625 ( .A(n28463), .B(img[584]), .S(n28581), .O(n12948) );
  AOI22S U30626 ( .A1(n28412), .A2(img[72]), .B1(n13775), .B2(n31714), .O(
        n28464) );
  ND2S U30627 ( .I1(n13808), .I2(n28464), .O(n28465) );
  MUX2 U30628 ( .A(img[48]), .B(n28465), .S(n28584), .O(n13484) );
  AOI22S U30629 ( .A1(n28347), .A2(img[48]), .B1(n24755), .B2(n31715), .O(
        n28466) );
  ND2S U30630 ( .I1(n13808), .I2(n28466), .O(n28467) );
  AOI22S U30631 ( .A1(n27065), .A2(img[968]), .B1(n13781), .B2(n31716), .O(
        n28469) );
  ND2S U30632 ( .I1(n13808), .I2(n28469), .O(n28470) );
  AOI22S U30633 ( .A1(n28106), .A2(img[944]), .B1(n24755), .B2(n31717), .O(
        n28471) );
  ND2S U30634 ( .I1(n13808), .I2(n28471), .O(n28472) );
  MUX2 U30635 ( .A(img[968]), .B(n28472), .S(n28623), .O(n12564) );
  AOI22S U30636 ( .A1(n27990), .A2(img[200]), .B1(n24755), .B2(n31718), .O(
        n28473) );
  ND2S U30637 ( .I1(n13808), .I2(n28473), .O(n28474) );
  MUX2 U30638 ( .A(img[176]), .B(n28474), .S(n28626), .O(n13356) );
  AOI22S U30639 ( .A1(n24415), .A2(img[176]), .B1(n24755), .B2(n31719), .O(
        n28475) );
  ND2S U30640 ( .I1(n13808), .I2(n28475), .O(n28476) );
  MUX2 U30641 ( .A(img[200]), .B(n28476), .S(n28629), .O(n13332) );
  AOI22S U30642 ( .A1(n26822), .A2(img[328]), .B1(n24755), .B2(n31720), .O(
        n28477) );
  ND2S U30643 ( .I1(n13808), .I2(n28477), .O(n28478) );
  MUX2 U30644 ( .A(img[304]), .B(n28478), .S(n28632), .O(n13228) );
  AOI22S U30645 ( .A1(n28083), .A2(img[304]), .B1(n25859), .B2(n31721), .O(
        n28479) );
  ND2S U30646 ( .I1(n28425), .I2(n28479), .O(n28480) );
  AOI22S U30647 ( .A1(n28347), .A2(img[456]), .B1(n25859), .B2(n31722), .O(
        n28481) );
  ND2S U30648 ( .I1(n28425), .I2(n28481), .O(n28482) );
  AOI22S U30649 ( .A1(n26970), .A2(img[432]), .B1(n29194), .B2(n31723), .O(
        n28483) );
  ND2S U30650 ( .I1(n28425), .I2(n28483), .O(n28484) );
  MUX2 U30651 ( .A(n28484), .B(img[456]), .S(n28641), .O(n13076) );
  AOI22S U30652 ( .A1(n26855), .A2(img[840]), .B1(n28433), .B2(n31724), .O(
        n28485) );
  ND2S U30653 ( .I1(n28425), .I2(n28485), .O(n28486) );
  INV1S U30654 ( .I(img[840]), .O(n28487) );
  AOI22S U30655 ( .A1(n29435), .A2(img[816]), .B1(n28162), .B2(n28487), .O(
        n28488) );
  ND2S U30656 ( .I1(n28425), .I2(n28488), .O(n28489) );
  AOI22S U30657 ( .A1(n24415), .A2(img[712]), .B1(n28862), .B2(n31725), .O(
        n28490) );
  ND2S U30658 ( .I1(n28425), .I2(n28490), .O(n28491) );
  AOI22S U30659 ( .A1(n28442), .A2(img[688]), .B1(n28913), .B2(n31726), .O(
        n28492) );
  ND2S U30660 ( .I1(n28425), .I2(n28492), .O(n28493) );
  AOI22S U30661 ( .A1(n29072), .A2(img[608]), .B1(n24755), .B2(n31727), .O(
        n28494) );
  ND2S U30662 ( .I1(n28425), .I2(n28494), .O(n28495) );
  AOI22S U30663 ( .A1(n26855), .A2(img[536]), .B1(n24193), .B2(n31728), .O(
        n28496) );
  ND2S U30664 ( .I1(n28292), .I2(n28496), .O(n28497) );
  AOI22S U30665 ( .A1(n28347), .A2(img[96]), .B1(n24193), .B2(n31729), .O(
        n28498) );
  ND2S U30666 ( .I1(n28425), .I2(n28498), .O(n28499) );
  AOI22S U30667 ( .A1(n13773), .A2(img[24]), .B1(n29407), .B2(n31730), .O(
        n28500) );
  ND2S U30668 ( .I1(n28425), .I2(n28500), .O(n28501) );
  MUX2 U30669 ( .A(img[96]), .B(n28501), .S(n29280), .O(n13436) );
  AOI22S U30670 ( .A1(n13777), .A2(img[992]), .B1(n24193), .B2(n31731), .O(
        n28502) );
  ND2S U30671 ( .I1(n28425), .I2(n28502), .O(n28503) );
  AOI22S U30672 ( .A1(n26970), .A2(img[920]), .B1(n23918), .B2(n31732), .O(
        n28504) );
  ND2S U30673 ( .I1(n28425), .I2(n28504), .O(n28505) );
  MUX2 U30674 ( .A(img[992]), .B(n28505), .S(n29224), .O(n12540) );
  AOI22S U30675 ( .A1(n28347), .A2(img[224]), .B1(n28913), .B2(n31733), .O(
        n28506) );
  ND2S U30676 ( .I1(n28425), .I2(n28506), .O(n28507) );
  MUX2 U30677 ( .A(img[152]), .B(n28507), .S(n29264), .O(n13380) );
  AOI22S U30678 ( .A1(n13777), .A2(img[152]), .B1(n23918), .B2(n31734), .O(
        n28508) );
  ND2S U30679 ( .I1(n28425), .I2(n28508), .O(n28509) );
  MUX2 U30680 ( .A(img[224]), .B(n28509), .S(n29267), .O(n13308) );
  AOI22S U30681 ( .A1(n13771), .A2(img[352]), .B1(n28862), .B2(n31735), .O(
        n28510) );
  ND2S U30682 ( .I1(n28425), .I2(n28510), .O(n28511) );
  AOI22S U30683 ( .A1(n13778), .A2(img[280]), .B1(n28862), .B2(n31736), .O(
        n28512) );
  ND2S U30684 ( .I1(n28425), .I2(n28512), .O(n28513) );
  MUX2 U30685 ( .A(img[352]), .B(n28513), .S(n29182), .O(n13180) );
  AOI22S U30686 ( .A1(n28318), .A2(img[480]), .B1(n24755), .B2(n31737), .O(
        n28514) );
  ND2S U30687 ( .I1(n28425), .I2(n28514), .O(n28515) );
  AOI22S U30688 ( .A1(n28382), .A2(img[408]), .B1(n28433), .B2(n31738), .O(
        n28516) );
  ND2S U30689 ( .I1(n28425), .I2(n28516), .O(n28517) );
  AOI22S U30690 ( .A1(n28643), .A2(img[864]), .B1(n13781), .B2(n31739), .O(
        n28518) );
  ND2S U30691 ( .I1(n28425), .I2(n28518), .O(n28519) );
  MUX2 U30692 ( .A(img[792]), .B(n28519), .S(n29227), .O(n12740) );
  INV1S U30693 ( .I(img[864]), .O(n28520) );
  AOI22S U30694 ( .A1(n28318), .A2(img[792]), .B1(n28862), .B2(n28520), .O(
        n28521) );
  ND2S U30695 ( .I1(n28425), .I2(n28521), .O(n28522) );
  AOI22S U30696 ( .A1(n29072), .A2(img[736]), .B1(n24755), .B2(n31740), .O(
        n28523) );
  ND2S U30697 ( .I1(n28425), .I2(n28523), .O(n28524) );
  AOI22S U30698 ( .A1(n29414), .A2(img[664]), .B1(n25062), .B2(n31741), .O(
        n28525) );
  ND2S U30699 ( .I1(n28425), .I2(n28525), .O(n28526) );
  OAI22S U30700 ( .A1(n28531), .A2(n28530), .B1(n13897), .B2(n28528), .O(
        n28532) );
  ND2S U30701 ( .I1(n28547), .I2(A67_shift[236]), .O(n28539) );
  AOI22S U30702 ( .A1(n28552), .A2(A67_shift[140]), .B1(n28551), .B2(
        A67_shift[204]), .O(n28538) );
  ND2S U30703 ( .I1(n28554), .I2(A67_shift[108]), .O(n28537) );
  INV1S U30704 ( .I(A67_shift[44]), .O(n28543) );
  AOI22S U30705 ( .A1(n28553), .A2(A67_shift[12]), .B1(n28546), .B2(
        A67_shift[172]), .O(n28542) );
  AOI12HS U30706 ( .B1(n28550), .B2(A67_shift[76]), .A1(n28540), .O(n28541) );
  OAI112HS U30707 ( .C1(n28544), .C2(n28543), .A1(n28542), .B1(n28541), .O(
        n28562) );
  AOI22S U30708 ( .A1(n28546), .A2(A67_shift[188]), .B1(n28545), .B2(
        A67_shift[60]), .O(n28549) );
  ND2S U30709 ( .I1(n28550), .I2(A67_shift[92]), .O(n28559) );
  AOI22S U30710 ( .A1(n28552), .A2(A67_shift[156]), .B1(n28551), .B2(
        A67_shift[220]), .O(n28558) );
  AOI22S U30711 ( .A1(n28554), .A2(A67_shift[124]), .B1(n28553), .B2(
        A67_shift[28]), .O(n28556) );
  AN2B1S U30712 ( .I1(n28556), .B1(n28555), .O(n28557) );
  OAI22S U30713 ( .A1(n28563), .A2(n28562), .B1(n28561), .B2(n28560), .O(
        n28572) );
  ND2S U30714 ( .I1(n28564), .I2(gray_avg_out[4]), .O(n28569) );
  ND2S U30715 ( .I1(n28565), .I2(gray_weight_out[4]), .O(n28568) );
  ND2S U30716 ( .I1(n28566), .I2(gray_max_out[4]), .O(n28567) );
  AOI22S U30717 ( .A1(n13778), .A2(img[588]), .B1(n23941), .B2(n31742), .O(
        n28577) );
  ND2S U30718 ( .I1(n29197), .I2(n28577), .O(n28579) );
  MUX2 U30719 ( .A(n28579), .B(img[564]), .S(n28578), .O(n12968) );
  AOI22S U30720 ( .A1(n28347), .A2(img[564]), .B1(n24374), .B2(n31743), .O(
        n28580) );
  ND2S U30721 ( .I1(n29197), .I2(n28580), .O(n28582) );
  MUX2 U30722 ( .A(n28582), .B(img[588]), .S(n28581), .O(n12944) );
  AOI22S U30723 ( .A1(n26855), .A2(img[76]), .B1(n13775), .B2(n31744), .O(
        n28583) );
  ND2S U30724 ( .I1(n29197), .I2(n28583), .O(n28585) );
  MUX2 U30725 ( .A(img[52]), .B(n28585), .S(n28584), .O(n13477) );
  AOI22S U30726 ( .A1(n29129), .A2(img[52]), .B1(n13775), .B2(n31745), .O(
        n28586) );
  ND2S U30727 ( .I1(n29197), .I2(n28586), .O(n28588) );
  MUX2 U30728 ( .A(img[76]), .B(n28588), .S(n28587), .O(n13456) );
  AOI22S U30729 ( .A1(n28347), .A2(img[1268]), .B1(n13775), .B2(n31746), .O(
        n28589) );
  ND2S U30730 ( .I1(n29197), .I2(n28589), .O(n28591) );
  MUX2 U30731 ( .A(img[1164]), .B(n28591), .S(n28590), .O(n12368) );
  AOI22S U30732 ( .A1(n28592), .A2(n31747), .B1(n27919), .B2(img[1164]), .O(
        n28594) );
  ND3S U30733 ( .I1(n29197), .I2(n28594), .I3(n28593), .O(n28596) );
  MUX2 U30734 ( .A(img[1268]), .B(n28596), .S(n28595), .O(n12264) );
  AOI22S U30735 ( .A1(n27990), .A2(img[1228]), .B1(n13775), .B2(n31748), .O(
        n28597) );
  ND2S U30736 ( .I1(n29197), .I2(n28597), .O(n28599) );
  AOI22S U30737 ( .A1(n29096), .A2(n31749), .B1(n28254), .B2(img[1204]), .O(
        n28601) );
  ND2S U30738 ( .I1(n29124), .I2(img[1268]), .O(n28600) );
  ND3S U30739 ( .I1(n29197), .I2(n28601), .I3(n28600), .O(n28603) );
  MUX2 U30740 ( .A(img[1228]), .B(n28603), .S(n28602), .O(n12304) );
  AOI22S U30741 ( .A1(n13771), .A2(img[1396]), .B1(n13775), .B2(n31750), .O(
        n28604) );
  ND2S U30742 ( .I1(n29197), .I2(n28604), .O(n28606) );
  MUX2 U30743 ( .A(img[1292]), .B(n28606), .S(n28605), .O(n12240) );
  AOI22S U30744 ( .A1(n28614), .A2(n31751), .B1(n27919), .B2(img[1292]), .O(
        n28608) );
  ND2S U30745 ( .I1(n13819), .I2(img[1356]), .O(n28607) );
  ND3S U30746 ( .I1(n29197), .I2(n28608), .I3(n28607), .O(n28610) );
  MUX2 U30747 ( .A(img[1396]), .B(n28610), .S(n28609), .O(n12136) );
  AOI22S U30748 ( .A1(n28347), .A2(img[1356]), .B1(n13775), .B2(n31752), .O(
        n28611) );
  ND2S U30749 ( .I1(n29197), .I2(n28611), .O(n28613) );
  MUX2 U30750 ( .A(n28613), .B(img[1332]), .S(n28612), .O(n12200) );
  AOI22S U30751 ( .A1(n28614), .A2(n31753), .B1(n24313), .B2(img[1332]), .O(
        n28616) );
  ND3S U30752 ( .I1(n29197), .I2(n28616), .I3(n28615), .O(n28618) );
  MUX2 U30753 ( .A(img[1356]), .B(n28618), .S(n28617), .O(n12176) );
  AOI22S U30754 ( .A1(n27065), .A2(img[972]), .B1(n13775), .B2(n31754), .O(
        n28619) );
  ND2S U30755 ( .I1(n29197), .I2(n28619), .O(n28621) );
  AOI22S U30756 ( .A1(n28643), .A2(img[948]), .B1(n25859), .B2(n31755), .O(
        n28622) );
  ND2S U30757 ( .I1(n29197), .I2(n28622), .O(n28624) );
  MUX2 U30758 ( .A(img[972]), .B(n28624), .S(n28623), .O(n12560) );
  AOI22S U30759 ( .A1(n28318), .A2(img[204]), .B1(n25591), .B2(n31756), .O(
        n28625) );
  ND2S U30760 ( .I1(n29197), .I2(n28625), .O(n28627) );
  MUX2 U30761 ( .A(img[180]), .B(n28627), .S(n28626), .O(n13352) );
  AOI22S U30762 ( .A1(n28318), .A2(img[180]), .B1(n25377), .B2(n31757), .O(
        n28628) );
  ND2S U30763 ( .I1(n29197), .I2(n28628), .O(n28630) );
  MUX2 U30764 ( .A(img[204]), .B(n28630), .S(n28629), .O(n13328) );
  AOI22S U30765 ( .A1(n28382), .A2(img[332]), .B1(n28433), .B2(n31758), .O(
        n28631) );
  ND2S U30766 ( .I1(n29197), .I2(n28631), .O(n28633) );
  MUX2 U30767 ( .A(img[308]), .B(n28633), .S(n28632), .O(n13224) );
  AOI22S U30768 ( .A1(n28382), .A2(img[308]), .B1(n13781), .B2(n31759), .O(
        n28634) );
  ND2S U30769 ( .I1(n29197), .I2(n28634), .O(n28636) );
  AOI22S U30770 ( .A1(n28382), .A2(img[460]), .B1(n25591), .B2(n31760), .O(
        n28637) );
  ND2S U30771 ( .I1(n29197), .I2(n28637), .O(n28639) );
  MUX2 U30772 ( .A(n28639), .B(img[436]), .S(n28638), .O(n13096) );
  AOI22S U30773 ( .A1(n28643), .A2(img[436]), .B1(n25062), .B2(n31761), .O(
        n28640) );
  ND2S U30774 ( .I1(n29197), .I2(n28640), .O(n28642) );
  AOI22S U30775 ( .A1(n28347), .A2(img[1524]), .B1(n28135), .B2(n31762), .O(
        n28644) );
  ND2S U30776 ( .I1(n29197), .I2(n28644), .O(n28646) );
  MUX2 U30777 ( .A(n28646), .B(img[1420]), .S(n28645), .O(n12112) );
  AOI22S U30778 ( .A1(n25591), .A2(n31763), .B1(n25444), .B2(img[1420]), .O(
        n28648) );
  ND3S U30779 ( .I1(n29197), .I2(n28648), .I3(n28647), .O(n28650) );
  AOI22S U30780 ( .A1(n27746), .A2(img[1484]), .B1(n13781), .B2(n31764), .O(
        n28651) );
  ND2S U30781 ( .I1(n29197), .I2(n28651), .O(n28653) );
  AOI22S U30782 ( .A1(n25591), .A2(n31765), .B1(n28043), .B2(img[1460]), .O(
        n28655) );
  ND2S U30783 ( .I1(n13820), .I2(img[1524]), .O(n28654) );
  AOI22S U30784 ( .A1(n26970), .A2(img[844]), .B1(n29194), .B2(n31766), .O(
        n28658) );
  ND2S U30785 ( .I1(n29197), .I2(n28658), .O(n28660) );
  INV1S U30786 ( .I(img[844]), .O(n28661) );
  AOI22S U30787 ( .A1(n28840), .A2(img[820]), .B1(n23918), .B2(n28661), .O(
        n28662) );
  ND2S U30788 ( .I1(n29197), .I2(n28662), .O(n28664) );
  MUX2 U30789 ( .A(n28664), .B(img[844]), .S(n28663), .O(n12688) );
  AOI22S U30790 ( .A1(n28347), .A2(img[716]), .B1(n28343), .B2(n31767), .O(
        n28665) );
  ND2S U30791 ( .I1(n29197), .I2(n28665), .O(n28667) );
  AOI22S U30792 ( .A1(n13771), .A2(img[692]), .B1(n28075), .B2(n31768), .O(
        n28668) );
  ND2S U30793 ( .I1(n29197), .I2(n28668), .O(n28670) );
  AOI22S U30794 ( .A1(n25595), .A2(img[1876]), .B1(n27511), .B2(n31769), .O(
        n28671) );
  ND2S U30795 ( .I1(n29197), .I2(n28671), .O(n28673) );
  MUX2 U30796 ( .A(n28673), .B(img[1836]), .S(n28672), .O(n11696) );
  AOI22S U30797 ( .A1(n24374), .A2(n31770), .B1(n28043), .B2(img[1836]), .O(
        n28675) );
  ND3S U30798 ( .I1(n29197), .I2(n28675), .I3(n28674), .O(n28677) );
  MUX2 U30799 ( .A(img[1876]), .B(n28677), .S(n28676), .O(n11656) );
  AOI22S U30800 ( .A1(n27990), .A2(img[1900]), .B1(n27511), .B2(n31771), .O(
        n28678) );
  ND2S U30801 ( .I1(n29197), .I2(n28678), .O(n28680) );
  MUX2 U30802 ( .A(n28680), .B(img[1812]), .S(n28679), .O(n11720) );
  AOI22S U30803 ( .A1(n28695), .A2(n31772), .B1(n28069), .B2(img[1812]), .O(
        n28682) );
  AOI22S U30804 ( .A1(n13770), .A2(img[1876]), .B1(img[1908]), .B2(n13782), 
        .O(n28681) );
  ND3S U30805 ( .I1(n29197), .I2(n28682), .I3(n28681), .O(n28684) );
  MUX2 U30806 ( .A(img[1900]), .B(n28684), .S(n28683), .O(n11632) );
  AOI22S U30807 ( .A1(n24415), .A2(img[1908]), .B1(n25062), .B2(n31773), .O(
        n28685) );
  ND2S U30808 ( .I1(n29197), .I2(n28685), .O(n28687) );
  AOI22S U30809 ( .A1(n28695), .A2(n31774), .B1(n25444), .B2(img[1804]), .O(
        n28689) );
  AOI22S U30810 ( .A1(n13819), .A2(img[1868]), .B1(img[1900]), .B2(n13782), 
        .O(n28688) );
  ND3S U30811 ( .I1(n29197), .I2(n28689), .I3(n28688), .O(n28691) );
  MUX2 U30812 ( .A(img[1908]), .B(n28691), .S(n28690), .O(n11624) );
  AOI22S U30813 ( .A1(n28840), .A2(img[1868]), .B1(n28592), .B2(n31775), .O(
        n28692) );
  ND2S U30814 ( .I1(n29197), .I2(n28692), .O(n28694) );
  MUX2 U30815 ( .A(n28694), .B(img[1844]), .S(n28693), .O(n11688) );
  AOI22S U30816 ( .A1(n28695), .A2(n31776), .B1(n25444), .B2(img[1844]), .O(
        n28697) );
  ND3S U30817 ( .I1(n29197), .I2(n28697), .I3(n28696), .O(n28699) );
  MUX2 U30818 ( .A(img[1868]), .B(n28699), .S(n28698), .O(n11664) );
  AOI22S U30819 ( .A1(n26822), .A2(img[1748]), .B1(n28695), .B2(n31777), .O(
        n28700) );
  ND2S U30820 ( .I1(n29197), .I2(n28700), .O(n28702) );
  AOI22S U30821 ( .A1(n29242), .A2(n31778), .B1(n25444), .B2(img[1708]), .O(
        n28704) );
  ND2S U30822 ( .I1(n29124), .I2(img[1772]), .O(n28703) );
  ND3S U30823 ( .I1(n29197), .I2(n28704), .I3(n28703), .O(n28706) );
  MUX2 U30824 ( .A(img[1748]), .B(n28706), .S(n28705), .O(n11784) );
  AOI22S U30825 ( .A1(n13778), .A2(img[1772]), .B1(n28592), .B2(n31779), .O(
        n28707) );
  ND2S U30826 ( .I1(n29197), .I2(n28707), .O(n28709) );
  MUX2 U30827 ( .A(n28709), .B(img[1684]), .S(n28708), .O(n11848) );
  AOI22S U30828 ( .A1(n29242), .A2(n31780), .B1(n25444), .B2(img[1684]), .O(
        n28711) );
  AOI22S U30829 ( .A1(n29124), .A2(img[1748]), .B1(img[1780]), .B2(n13782), 
        .O(n28710) );
  ND3S U30830 ( .I1(n29197), .I2(n28711), .I3(n28710), .O(n28713) );
  MUX2 U30831 ( .A(img[1772]), .B(n28713), .S(n28712), .O(n11760) );
  AOI22S U30832 ( .A1(n24415), .A2(img[1780]), .B1(n28135), .B2(n31781), .O(
        n28714) );
  ND2S U30833 ( .I1(n29197), .I2(n28714), .O(n28716) );
  MUX2 U30834 ( .A(img[1676]), .B(n28716), .S(n28715), .O(n11856) );
  AOI22S U30835 ( .A1(n25591), .A2(n31782), .B1(n25444), .B2(img[1676]), .O(
        n28718) );
  AOI22S U30836 ( .A1(n13905), .A2(img[1740]), .B1(img[1772]), .B2(n13782), 
        .O(n28717) );
  ND3S U30837 ( .I1(n29197), .I2(n28718), .I3(n28717), .O(n28720) );
  MUX2 U30838 ( .A(img[1780]), .B(n28720), .S(n28719), .O(n11752) );
  AOI22S U30839 ( .A1(n27746), .A2(img[1740]), .B1(n29530), .B2(n31783), .O(
        n28721) );
  ND2S U30840 ( .I1(n29197), .I2(n28721), .O(n28723) );
  MUX2 U30841 ( .A(n28723), .B(img[1716]), .S(n28722), .O(n11816) );
  AOI22S U30842 ( .A1(n29242), .A2(n31784), .B1(n25444), .B2(img[1716]), .O(
        n28725) );
  ND2S U30843 ( .I1(n13770), .I2(img[1780]), .O(n28724) );
  ND3S U30844 ( .I1(n29197), .I2(n28725), .I3(n28724), .O(n28727) );
  MUX2 U30845 ( .A(img[1740]), .B(n28727), .S(n28726), .O(n11792) );
  AOI22S U30846 ( .A1(n25595), .A2(img[1620]), .B1(n28182), .B2(n31785), .O(
        n28728) );
  ND2S U30847 ( .I1(n29197), .I2(n28728), .O(n28730) );
  MUX2 U30848 ( .A(n28730), .B(img[1580]), .S(n28729), .O(n11952) );
  AOI22S U30849 ( .A1(n13779), .A2(n31786), .B1(n28069), .B2(img[1580]), .O(
        n28732) );
  ND2S U30850 ( .I1(n13819), .I2(img[1644]), .O(n28731) );
  ND3S U30851 ( .I1(n29197), .I2(n28732), .I3(n28731), .O(n28734) );
  MUX2 U30852 ( .A(img[1620]), .B(n28734), .S(n28733), .O(n11912) );
  AOI22S U30853 ( .A1(n28347), .A2(img[1644]), .B1(n25062), .B2(n31787), .O(
        n28735) );
  ND2S U30854 ( .I1(n29197), .I2(n28735), .O(n28737) );
  MUX2 U30855 ( .A(n28737), .B(img[1556]), .S(n28736), .O(n11976) );
  BUF12CK U30856 ( .I(n29278), .O(n29197) );
  AOI22S U30857 ( .A1(n29530), .A2(n31788), .B1(n24946), .B2(img[1556]), .O(
        n28739) );
  AOI22S U30858 ( .A1(n13902), .A2(img[1620]), .B1(img[1652]), .B2(n13782), 
        .O(n28738) );
  ND3S U30859 ( .I1(n29197), .I2(n28739), .I3(n28738), .O(n28741) );
  MUX2 U30860 ( .A(img[1644]), .B(n28741), .S(n28740), .O(n11888) );
  AOI22S U30861 ( .A1(n26101), .A2(img[1652]), .B1(n24755), .B2(n31789), .O(
        n28742) );
  ND2S U30862 ( .I1(n29197), .I2(n28742), .O(n28744) );
  AOI22S U30863 ( .A1(n28162), .A2(n31790), .B1(n28254), .B2(img[1548]), .O(
        n28746) );
  AOI22S U30864 ( .A1(n13903), .A2(img[1612]), .B1(img[1644]), .B2(n13782), 
        .O(n28745) );
  ND3S U30865 ( .I1(n29197), .I2(n28746), .I3(n28745), .O(n28748) );
  MUX2 U30866 ( .A(img[1652]), .B(n28748), .S(n28747), .O(n11880) );
  AOI22S U30867 ( .A1(n13777), .A2(img[1612]), .B1(n28695), .B2(n31791), .O(
        n28749) );
  ND2S U30868 ( .I1(n29197), .I2(n28749), .O(n28751) );
  AOI22S U30869 ( .A1(n29457), .A2(n31792), .B1(n24313), .B2(img[1588]), .O(
        n28753) );
  ND2S U30870 ( .I1(n29124), .I2(img[1652]), .O(n28752) );
  ND3S U30871 ( .I1(n29197), .I2(n28753), .I3(n28752), .O(n28755) );
  MUX2 U30872 ( .A(img[1612]), .B(n28755), .S(n28754), .O(n11920) );
  AOI22S U30873 ( .A1(n27065), .A2(img[1140]), .B1(n29096), .B2(n31793), .O(
        n28756) );
  ND2S U30874 ( .I1(n29197), .I2(n28756), .O(n28758) );
  MUX2 U30875 ( .A(img[1036]), .B(n28758), .S(n28757), .O(n12496) );
  AOI22S U30876 ( .A1(n27735), .A2(n31794), .B1(n25444), .B2(img[1036]), .O(
        n28760) );
  ND2S U30877 ( .I1(n13770), .I2(img[1100]), .O(n28759) );
  ND3S U30878 ( .I1(n29197), .I2(n28760), .I3(n28759), .O(n28762) );
  MUX2 U30879 ( .A(img[1140]), .B(n28762), .S(n28761), .O(n12392) );
  AOI22S U30880 ( .A1(n13780), .A2(img[1100]), .B1(n29194), .B2(n31795), .O(
        n28763) );
  ND2S U30881 ( .I1(n29197), .I2(n28763), .O(n28765) );
  MUX2 U30882 ( .A(n28765), .B(img[1076]), .S(n28764), .O(n12456) );
  AOI22S U30883 ( .A1(n27735), .A2(n31796), .B1(n24946), .B2(img[1076]), .O(
        n28767) );
  ND3S U30884 ( .I1(n29197), .I2(n28767), .I3(n28766), .O(n28769) );
  MUX2 U30885 ( .A(img[1100]), .B(n28769), .S(n28768), .O(n12432) );
  AOI22S U30886 ( .A1(n28840), .A2(img[2004]), .B1(n28862), .B2(n31797), .O(
        n28770) );
  ND2S U30887 ( .I1(n29197), .I2(n28770), .O(n28772) );
  AOI22S U30888 ( .A1(n28433), .A2(n31798), .B1(n28254), .B2(img[1964]), .O(
        n28774) );
  ND2S U30889 ( .I1(n13820), .I2(img[2028]), .O(n28773) );
  ND3S U30890 ( .I1(n29197), .I2(n28774), .I3(n28773), .O(n28776) );
  MUX2 U30891 ( .A(img[2004]), .B(n28776), .S(n28775), .O(n11528) );
  AOI22S U30892 ( .A1(n13772), .A2(img[2028]), .B1(n25062), .B2(n31799), .O(
        n28777) );
  ND2S U30893 ( .I1(n29197), .I2(n28777), .O(n28779) );
  MUX2 U30894 ( .A(n28779), .B(img[1940]), .S(n28778), .O(n11592) );
  AOI22S U30895 ( .A1(n28135), .A2(n31800), .B1(n24313), .B2(img[1940]), .O(
        n28781) );
  AOI22S U30896 ( .A1(n13899), .A2(img[2004]), .B1(img[2036]), .B2(n13782), 
        .O(n28780) );
  ND3S U30897 ( .I1(n29197), .I2(n28781), .I3(n28780), .O(n28783) );
  MUX2 U30898 ( .A(img[2028]), .B(n28783), .S(n28782), .O(n11504) );
  AOI22S U30899 ( .A1(n26855), .A2(img[2036]), .B1(n28135), .B2(n31801), .O(
        n28784) );
  ND2S U30900 ( .I1(n29197), .I2(n28784), .O(n28786) );
  MUX2 U30901 ( .A(img[1932]), .B(n28786), .S(n28785), .O(n11600) );
  AOI22S U30902 ( .A1(n28695), .A2(n31802), .B1(n27919), .B2(img[1932]), .O(
        n28788) );
  AOI22S U30903 ( .A1(n13903), .A2(img[1996]), .B1(img[2028]), .B2(n13782), 
        .O(n28787) );
  ND3S U30904 ( .I1(n29197), .I2(n28788), .I3(n28787), .O(n28790) );
  MUX2 U30905 ( .A(img[2036]), .B(n28790), .S(n28789), .O(n11496) );
  AOI22S U30906 ( .A1(n29072), .A2(img[1996]), .B1(n27511), .B2(n31803), .O(
        n28791) );
  ND2S U30907 ( .I1(n29197), .I2(n28791), .O(n28793) );
  MUX2 U30908 ( .A(n28793), .B(img[1972]), .S(n28792), .O(n11560) );
  AOI22S U30909 ( .A1(n29096), .A2(n31804), .B1(n28069), .B2(img[1972]), .O(
        n28795) );
  ND3S U30910 ( .I1(n29197), .I2(n28795), .I3(n28794), .O(n28797) );
  MUX2 U30911 ( .A(img[1996]), .B(n28797), .S(n28796), .O(n11536) );
  AOI22S U30912 ( .A1(n26101), .A2(img[572]), .B1(n28592), .B2(n31805), .O(
        n28798) );
  ND2S U30913 ( .I1(n29197), .I2(n28798), .O(n28800) );
  MUX2 U30914 ( .A(n28800), .B(img[580]), .S(n28799), .O(n12952) );
  AOI22S U30915 ( .A1(n28083), .A2(img[580]), .B1(n28592), .B2(n31806), .O(
        n28801) );
  ND2S U30916 ( .I1(n29197), .I2(n28801), .O(n28802) );
  MUX2 U30917 ( .A(n28802), .B(img[572]), .S(n29532), .O(n12960) );
  AOI22S U30918 ( .A1(n25595), .A2(img[60]), .B1(n27511), .B2(n31807), .O(
        n28803) );
  ND2S U30919 ( .I1(n29197), .I2(n28803), .O(n28805) );
  MUX2 U30920 ( .A(img[68]), .B(n28805), .S(n28804), .O(n13464) );
  AOI22S U30921 ( .A1(n28106), .A2(img[68]), .B1(n28592), .B2(n31808), .O(
        n28806) );
  ND2S U30922 ( .I1(n29197), .I2(n28806), .O(n28808) );
  MUX2 U30923 ( .A(img[60]), .B(n28808), .S(n28807), .O(n13472) );
  AOI22S U30924 ( .A1(n26101), .A2(img[1276]), .B1(n28862), .B2(n31809), .O(
        n28809) );
  ND2S U30925 ( .I1(n29197), .I2(n28809), .O(n28811) );
  MUX2 U30926 ( .A(img[1156]), .B(n28811), .S(n28810), .O(n12376) );
  AOI22S U30927 ( .A1(n13781), .A2(n31810), .B1(n25444), .B2(img[1156]), .O(
        n28813) );
  ND3S U30928 ( .I1(n29197), .I2(n28813), .I3(n28812), .O(n28815) );
  MUX2 U30929 ( .A(img[1276]), .B(n28815), .S(n28814), .O(n12256) );
  AOI22S U30930 ( .A1(n28913), .A2(n31811), .B1(n27919), .B2(img[1212]), .O(
        n28817) );
  ND2S U30931 ( .I1(n13770), .I2(img[1276]), .O(n28816) );
  ND3S U30932 ( .I1(n29197), .I2(n28817), .I3(n28816), .O(n28819) );
  MUX2 U30933 ( .A(img[1220]), .B(n28819), .S(n28818), .O(n12312) );
  AOI22S U30934 ( .A1(n28840), .A2(img[1220]), .B1(n29397), .B2(n31812), .O(
        n28820) );
  ND2S U30935 ( .I1(n29197), .I2(n28820), .O(n28822) );
  MUX2 U30936 ( .A(img[1212]), .B(n28822), .S(n28821), .O(n12320) );
  AOI22S U30937 ( .A1(n13780), .A2(img[1404]), .B1(n28614), .B2(n31813), .O(
        n28823) );
  ND2S U30938 ( .I1(n29197), .I2(n28823), .O(n28825) );
  MUX2 U30939 ( .A(img[1284]), .B(n28825), .S(n28824), .O(n12248) );
  AOI22S U30940 ( .A1(n28913), .A2(n31814), .B1(n24313), .B2(img[1284]), .O(
        n28827) );
  ND3S U30941 ( .I1(n29197), .I2(n28827), .I3(n28826), .O(n28829) );
  MUX2 U30942 ( .A(img[1404]), .B(n28829), .S(n28828), .O(n12128) );
  AOI22S U30943 ( .A1(n25062), .A2(n31815), .B1(n25444), .B2(img[1340]), .O(
        n28831) );
  ND3S U30944 ( .I1(n29197), .I2(n28831), .I3(n28830), .O(n28833) );
  MUX2 U30945 ( .A(img[1348]), .B(n28833), .S(n28832), .O(n12184) );
  AOI22S U30946 ( .A1(n13776), .A2(img[1348]), .B1(n29194), .B2(n31816), .O(
        n28834) );
  ND2S U30947 ( .I1(n29197), .I2(n28834), .O(n28836) );
  AOI22S U30948 ( .A1(n28106), .A2(img[956]), .B1(n13781), .B2(n31817), .O(
        n28837) );
  ND2S U30949 ( .I1(n29197), .I2(n28837), .O(n28839) );
  MUX2 U30950 ( .A(img[964]), .B(n28839), .S(n28838), .O(n12568) );
  AOI22S U30951 ( .A1(n28840), .A2(img[964]), .B1(n25062), .B2(n31818), .O(
        n28841) );
  ND2S U30952 ( .I1(n29197), .I2(n28841), .O(n28843) );
  AOI22S U30953 ( .A1(n28840), .A2(img[188]), .B1(n13779), .B2(n31819), .O(
        n28844) );
  ND2S U30954 ( .I1(n29197), .I2(n28844), .O(n28846) );
  MUX2 U30955 ( .A(img[196]), .B(n28846), .S(n28845), .O(n13336) );
  AOI22S U30956 ( .A1(n28840), .A2(img[196]), .B1(n28433), .B2(n31820), .O(
        n28847) );
  ND2S U30957 ( .I1(n29197), .I2(n28847), .O(n28849) );
  MUX2 U30958 ( .A(img[188]), .B(n28849), .S(n28848), .O(n13344) );
  AOI22S U30959 ( .A1(n28840), .A2(img[316]), .B1(n13781), .B2(n31821), .O(
        n28850) );
  ND2S U30960 ( .I1(n29197), .I2(n28850), .O(n28852) );
  MUX2 U30961 ( .A(img[324]), .B(n28852), .S(n28851), .O(n13208) );
  AOI22S U30962 ( .A1(n26822), .A2(img[324]), .B1(n28913), .B2(n31822), .O(
        n28853) );
  ND2S U30963 ( .I1(n29197), .I2(n28853), .O(n28855) );
  AOI22S U30964 ( .A1(n26822), .A2(img[444]), .B1(n25591), .B2(n31823), .O(
        n28856) );
  ND2S U30965 ( .I1(n13806), .I2(n28856), .O(n28858) );
  MUX2 U30966 ( .A(img[452]), .B(n28858), .S(n28857), .O(n13080) );
  AOI22S U30967 ( .A1(n26101), .A2(img[452]), .B1(n29242), .B2(n31824), .O(
        n28859) );
  ND2S U30968 ( .I1(n13806), .I2(n28859), .O(n28861) );
  MUX2 U30969 ( .A(img[444]), .B(n28861), .S(n28860), .O(n13089) );
  AOI22S U30970 ( .A1(n28347), .A2(img[1532]), .B1(n28433), .B2(n31825), .O(
        n28863) );
  ND2S U30971 ( .I1(n13806), .I2(n28863), .O(n28865) );
  MUX2 U30972 ( .A(img[1412]), .B(n28865), .S(n28864), .O(n12120) );
  AOI22S U30973 ( .A1(n24374), .A2(n31826), .B1(n28254), .B2(img[1412]), .O(
        n28867) );
  ND2S U30974 ( .I1(n13770), .I2(img[1476]), .O(n28866) );
  ND3S U30975 ( .I1(n29197), .I2(n28867), .I3(n28866), .O(n28869) );
  AOI22S U30976 ( .A1(n28182), .A2(n31827), .B1(n24313), .B2(img[1468]), .O(
        n28871) );
  ND2S U30977 ( .I1(n29124), .I2(img[1532]), .O(n28870) );
  ND3S U30978 ( .I1(n29197), .I2(n28871), .I3(n28870), .O(n28873) );
  MUX2 U30979 ( .A(img[1476]), .B(n28873), .S(n28872), .O(n12056) );
  AOI22S U30980 ( .A1(n13773), .A2(img[1476]), .B1(n25591), .B2(n31828), .O(
        n28874) );
  ND2S U30981 ( .I1(n13806), .I2(n28874), .O(n28876) );
  INV1S U30982 ( .I(img[836]), .O(n28877) );
  AOI22S U30983 ( .A1(n29435), .A2(img[828]), .B1(n27735), .B2(n28877), .O(
        n28878) );
  ND2S U30984 ( .I1(n13806), .I2(n28878), .O(n28880) );
  MUX2 U30985 ( .A(n28880), .B(img[836]), .S(n28879), .O(n12696) );
  INV1S U30986 ( .I(img[828]), .O(n28881) );
  AOI22S U30987 ( .A1(n28382), .A2(img[836]), .B1(n28862), .B2(n28881), .O(
        n28882) );
  ND2S U30988 ( .I1(n13806), .I2(n28882), .O(n28884) );
  AOI22S U30989 ( .A1(n13771), .A2(img[700]), .B1(n28862), .B2(n31829), .O(
        n28885) );
  ND2S U30990 ( .I1(n13806), .I2(n28885), .O(n28887) );
  AOI22S U30991 ( .A1(n13771), .A2(img[708]), .B1(n28862), .B2(n31830), .O(
        n28888) );
  ND2S U30992 ( .I1(n13806), .I2(n28888), .O(n28890) );
  AOI22S U30993 ( .A1(n13771), .A2(img[1884]), .B1(n28862), .B2(n31831), .O(
        n28891) );
  ND2S U30994 ( .I1(n13806), .I2(n28891), .O(n28893) );
  MUX2 U30995 ( .A(n28893), .B(img[1828]), .S(n28892), .O(n11704) );
  AOI22S U30996 ( .A1(n25377), .A2(n31832), .B1(n28069), .B2(img[1828]), .O(
        n28895) );
  ND2S U30997 ( .I1(n13819), .I2(img[1892]), .O(n28894) );
  ND3S U30998 ( .I1(n29197), .I2(n28895), .I3(n28894), .O(n28897) );
  AOI22S U30999 ( .A1(n13771), .A2(img[1892]), .B1(n28862), .B2(n31833), .O(
        n28898) );
  ND2S U31000 ( .I1(n13806), .I2(n28898), .O(n28900) );
  MUX2 U31001 ( .A(img[1820]), .B(n28900), .S(n28899), .O(n11712) );
  AOI22S U31002 ( .A1(n29194), .A2(n31834), .B1(n28043), .B2(img[1820]), .O(
        n28902) );
  AOI22S U31003 ( .A1(n13819), .A2(img[1884]), .B1(img[1916]), .B2(n13782), 
        .O(n28901) );
  ND3S U31004 ( .I1(n29197), .I2(n28902), .I3(n28901), .O(n28904) );
  MUX2 U31005 ( .A(img[1892]), .B(n28904), .S(n28903), .O(n11640) );
  AOI22S U31006 ( .A1(n28840), .A2(img[1916]), .B1(n28862), .B2(n31835), .O(
        n28905) );
  ND2S U31007 ( .I1(n13806), .I2(n28905), .O(n28907) );
  AOI22S U31008 ( .A1(n13779), .A2(n31836), .B1(n24313), .B2(img[1796]), .O(
        n28910) );
  AOI22S U31009 ( .A1(n29124), .A2(img[1860]), .B1(img[1892]), .B2(n28908), 
        .O(n28909) );
  ND3S U31010 ( .I1(n29197), .I2(n28910), .I3(n28909), .O(n28912) );
  MUX2 U31011 ( .A(img[1916]), .B(n28912), .S(n28911), .O(n11616) );
  AOI22S U31012 ( .A1(n28913), .A2(n31837), .B1(n28254), .B2(img[1852]), .O(
        n28915) );
  ND2S U31013 ( .I1(n13819), .I2(img[1916]), .O(n28914) );
  ND3S U31014 ( .I1(n29197), .I2(n28915), .I3(n28914), .O(n28917) );
  MUX2 U31015 ( .A(img[1860]), .B(n28917), .S(n28916), .O(n11672) );
  AOI22S U31016 ( .A1(n28840), .A2(img[1860]), .B1(n28862), .B2(n31838), .O(
        n28918) );
  ND2S U31017 ( .I1(n13806), .I2(n28918), .O(n28920) );
  MUX2 U31018 ( .A(img[1852]), .B(n28920), .S(n28919), .O(n11680) );
  AOI22S U31019 ( .A1(n28840), .A2(img[1756]), .B1(n28862), .B2(n31839), .O(
        n28921) );
  ND2S U31020 ( .I1(n13806), .I2(n28921), .O(n28923) );
  MUX2 U31021 ( .A(n28923), .B(img[1700]), .S(n28922), .O(n11832) );
  AOI22S U31022 ( .A1(n28135), .A2(n31840), .B1(n28069), .B2(img[1700]), .O(
        n28925) );
  ND2S U31023 ( .I1(n13770), .I2(img[1764]), .O(n28924) );
  ND3S U31024 ( .I1(n29197), .I2(n28925), .I3(n28924), .O(n28927) );
  AOI22S U31025 ( .A1(n28840), .A2(img[1764]), .B1(n28862), .B2(n31841), .O(
        n28928) );
  ND2S U31026 ( .I1(n13806), .I2(n28928), .O(n28930) );
  MUX2 U31027 ( .A(img[1692]), .B(n28930), .S(n28929), .O(n11840) );
  AOI22S U31028 ( .A1(n28614), .A2(n31842), .B1(n24946), .B2(img[1692]), .O(
        n28932) );
  AOI22S U31029 ( .A1(n29124), .A2(img[1756]), .B1(img[1788]), .B2(n13782), 
        .O(n28931) );
  ND3S U31030 ( .I1(n29197), .I2(n28932), .I3(n28931), .O(n28934) );
  MUX2 U31031 ( .A(img[1764]), .B(n28934), .S(n28933), .O(n11768) );
  AOI22S U31032 ( .A1(n28840), .A2(img[1788]), .B1(n29530), .B2(n31843), .O(
        n28935) );
  ND2S U31033 ( .I1(n13806), .I2(n28935), .O(n28937) );
  AOI22S U31034 ( .A1(n28938), .A2(n31844), .B1(n28069), .B2(img[1668]), .O(
        n28940) );
  AOI22S U31035 ( .A1(n13905), .A2(img[1732]), .B1(img[1764]), .B2(n13782), 
        .O(n28939) );
  ND3S U31036 ( .I1(n29197), .I2(n28940), .I3(n28939), .O(n28942) );
  MUX2 U31037 ( .A(img[1788]), .B(n28942), .S(n28941), .O(n11744) );
  AOI22S U31038 ( .A1(n13781), .A2(n31845), .B1(n28043), .B2(img[1724]), .O(
        n28944) );
  ND3S U31039 ( .I1(n29197), .I2(n28944), .I3(n28943), .O(n28946) );
  MUX2 U31040 ( .A(img[1732]), .B(n28946), .S(n28945), .O(n11800) );
  AOI22S U31041 ( .A1(n28840), .A2(img[1732]), .B1(n24755), .B2(n31846), .O(
        n28947) );
  ND2S U31042 ( .I1(n13806), .I2(n28947), .O(n28949) );
  MUX2 U31043 ( .A(img[1724]), .B(n28949), .S(n28948), .O(n11808) );
  AOI22S U31044 ( .A1(n28840), .A2(img[1628]), .B1(n24755), .B2(n31847), .O(
        n28950) );
  ND2S U31045 ( .I1(n13806), .I2(n28950), .O(n28952) );
  MUX2 U31046 ( .A(n28952), .B(img[1572]), .S(n28951), .O(n11960) );
  AOI22S U31047 ( .A1(n25468), .A2(n31848), .B1(n28069), .B2(img[1572]), .O(
        n28954) );
  ND2S U31048 ( .I1(n13819), .I2(img[1636]), .O(n28953) );
  ND3S U31049 ( .I1(n29197), .I2(n28954), .I3(n28953), .O(n28956) );
  BUF1 U31050 ( .I(n28318), .O(n29072) );
  AOI22S U31051 ( .A1(n29072), .A2(img[1636]), .B1(n24755), .B2(n31849), .O(
        n28957) );
  ND2S U31052 ( .I1(n13806), .I2(n28957), .O(n28959) );
  MUX2 U31053 ( .A(img[1564]), .B(n28959), .S(n28958), .O(n11968) );
  AOI22S U31054 ( .A1(n25591), .A2(n31850), .B1(n28069), .B2(img[1564]), .O(
        n28961) );
  AOI22S U31055 ( .A1(n29124), .A2(img[1628]), .B1(img[1660]), .B2(n13782), 
        .O(n28960) );
  ND3S U31056 ( .I1(n29197), .I2(n28961), .I3(n28960), .O(n28963) );
  MUX2 U31057 ( .A(img[1636]), .B(n28963), .S(n28962), .O(n11895) );
  AOI22S U31058 ( .A1(n29072), .A2(img[1660]), .B1(n28862), .B2(n31851), .O(
        n28964) );
  ND2S U31059 ( .I1(n13806), .I2(n28964), .O(n28966) );
  AOI22S U31060 ( .A1(n28075), .A2(n31852), .B1(n24313), .B2(img[1540]), .O(
        n28968) );
  AOI22S U31061 ( .A1(n13770), .A2(img[1604]), .B1(img[1636]), .B2(n13782), 
        .O(n28967) );
  ND3S U31062 ( .I1(n29197), .I2(n28968), .I3(n28967), .O(n28970) );
  MUX2 U31063 ( .A(img[1660]), .B(n28970), .S(n28969), .O(n11872) );
  AOI22S U31064 ( .A1(n28037), .A2(n31853), .B1(n24313), .B2(img[1596]), .O(
        n28972) );
  ND3S U31065 ( .I1(n29197), .I2(n28972), .I3(n28971), .O(n28974) );
  MUX2 U31066 ( .A(img[1604]), .B(n28974), .S(n28973), .O(n11928) );
  AOI22S U31067 ( .A1(n29072), .A2(img[1604]), .B1(n28913), .B2(n31854), .O(
        n28975) );
  ND2S U31068 ( .I1(n13806), .I2(n28975), .O(n28977) );
  MUX2 U31069 ( .A(img[1596]), .B(n28977), .S(n28976), .O(n11936) );
  AOI22S U31070 ( .A1(n29072), .A2(img[1148]), .B1(n25859), .B2(n31855), .O(
        n28978) );
  ND2S U31071 ( .I1(n13806), .I2(n28978), .O(n28980) );
  AOI22S U31072 ( .A1(n28135), .A2(n31856), .B1(n28069), .B2(img[1028]), .O(
        n28982) );
  ND2S U31073 ( .I1(n29124), .I2(img[1092]), .O(n28981) );
  ND3S U31074 ( .I1(n29197), .I2(n28982), .I3(n28981), .O(n28984) );
  MUX2 U31075 ( .A(img[1148]), .B(n28984), .S(n28983), .O(n12384) );
  AOI22S U31076 ( .A1(n28938), .A2(n31857), .B1(n24946), .B2(img[1084]), .O(
        n28986) );
  ND2S U31077 ( .I1(n13820), .I2(img[1148]), .O(n28985) );
  ND3S U31078 ( .I1(n29197), .I2(n28986), .I3(n28985), .O(n28988) );
  MUX2 U31079 ( .A(img[1092]), .B(n28988), .S(n28987), .O(n12437) );
  AOI22S U31080 ( .A1(n13771), .A2(img[1092]), .B1(n25468), .B2(n31858), .O(
        n28989) );
  ND2S U31081 ( .I1(n13806), .I2(n28989), .O(n28991) );
  AOI22S U31082 ( .A1(n13771), .A2(img[2012]), .B1(n13781), .B2(n31859), .O(
        n28992) );
  ND2S U31083 ( .I1(n13806), .I2(n28992), .O(n28994) );
  MUX2 U31084 ( .A(n28994), .B(img[1956]), .S(n28993), .O(n11576) );
  AOI22S U31085 ( .A1(n29194), .A2(n31860), .B1(n28254), .B2(img[1956]), .O(
        n28996) );
  ND3S U31086 ( .I1(n29197), .I2(n28996), .I3(n28995), .O(n28998) );
  AOI22S U31087 ( .A1(n13771), .A2(img[2020]), .B1(n29242), .B2(n31861), .O(
        n28999) );
  ND2S U31088 ( .I1(n13806), .I2(n28999), .O(n29001) );
  MUX2 U31089 ( .A(img[1948]), .B(n29001), .S(n29000), .O(n11584) );
  AOI22S U31090 ( .A1(n25591), .A2(n31862), .B1(n24946), .B2(img[1948]), .O(
        n29003) );
  AOI22S U31091 ( .A1(n29124), .A2(img[2012]), .B1(img[2044]), .B2(n13782), 
        .O(n29002) );
  ND3S U31092 ( .I1(n29197), .I2(n29003), .I3(n29002), .O(n29005) );
  MUX2 U31093 ( .A(img[2020]), .B(n29005), .S(n29004), .O(n11512) );
  AOI22S U31094 ( .A1(n13771), .A2(img[2044]), .B1(n28695), .B2(n31863), .O(
        n29006) );
  ND2S U31095 ( .I1(n13806), .I2(n29006), .O(n29008) );
  MUX2 U31096 ( .A(img[1924]), .B(n29008), .S(n29007), .O(n11608) );
  AOI22S U31097 ( .A1(n13779), .A2(n31864), .B1(n24946), .B2(img[1924]), .O(
        n29010) );
  AOI22S U31098 ( .A1(n13904), .A2(img[1988]), .B1(img[2020]), .B2(n13782), 
        .O(n29009) );
  ND3S U31099 ( .I1(n29197), .I2(n29010), .I3(n29009), .O(n29012) );
  AOI22S U31100 ( .A1(n28343), .A2(n31865), .B1(n29257), .B2(img[1980]), .O(
        n29014) );
  ND2S U31101 ( .I1(n13770), .I2(img[2044]), .O(n29013) );
  AOI22S U31102 ( .A1(n13771), .A2(img[1988]), .B1(n28913), .B2(n31866), .O(
        n29017) );
  ND2S U31103 ( .I1(n13806), .I2(n29017), .O(n29019) );
  MUX2 U31104 ( .A(img[1980]), .B(n29019), .S(n29018), .O(n11552) );
  AOI22S U31105 ( .A1(n13771), .A2(img[620]), .B1(n28614), .B2(n31867), .O(
        n29020) );
  ND2S U31106 ( .I1(n13806), .I2(n29020), .O(n29022) );
  AOI22S U31107 ( .A1(n13771), .A2(img[532]), .B1(n28913), .B2(n31868), .O(
        n29023) );
  ND2S U31108 ( .I1(n13806), .I2(n29023), .O(n29025) );
  MUX2 U31109 ( .A(n29025), .B(img[620]), .S(n29024), .O(n12912) );
  AOI22S U31110 ( .A1(n27990), .A2(img[108]), .B1(n25591), .B2(n31869), .O(
        n29026) );
  ND2S U31111 ( .I1(n13806), .I2(n29026), .O(n29028) );
  AOI22S U31112 ( .A1(n28318), .A2(img[20]), .B1(n27735), .B2(n31870), .O(
        n29029) );
  ND2S U31113 ( .I1(n13806), .I2(n29029), .O(n29031) );
  MUX2 U31114 ( .A(img[108]), .B(n29031), .S(n29030), .O(n13424) );
  AOI22S U31115 ( .A1(n28318), .A2(img[1236]), .B1(n29457), .B2(n31871), .O(
        n29032) );
  ND2S U31116 ( .I1(n13806), .I2(n29032), .O(n29034) );
  MUX2 U31117 ( .A(img[1196]), .B(n29034), .S(n29033), .O(n12336) );
  AOI22S U31118 ( .A1(n28037), .A2(n31872), .B1(n29257), .B2(img[1196]), .O(
        n29036) );
  ND3S U31119 ( .I1(n29197), .I2(n29036), .I3(n29035), .O(n29038) );
  MUX2 U31120 ( .A(img[1236]), .B(n29038), .S(n29037), .O(n12296) );
  AOI22S U31121 ( .A1(n28318), .A2(img[1260]), .B1(n13775), .B2(n31873), .O(
        n29039) );
  ND2S U31122 ( .I1(n13806), .I2(n29039), .O(n29041) );
  AOI22S U31123 ( .A1(n29096), .A2(n31874), .B1(n29257), .B2(img[1172]), .O(
        n29043) );
  ND2S U31124 ( .I1(n29124), .I2(img[1236]), .O(n29042) );
  ND3S U31125 ( .I1(n29197), .I2(n29043), .I3(n29042), .O(n29045) );
  MUX2 U31126 ( .A(img[1260]), .B(n29045), .S(n29044), .O(n12272) );
  AOI22S U31127 ( .A1(n29072), .A2(img[1364]), .B1(n25591), .B2(n31875), .O(
        n29046) );
  ND2S U31128 ( .I1(n13806), .I2(n29046), .O(n29048) );
  AOI22S U31129 ( .A1(n13779), .A2(n31876), .B1(n29257), .B2(img[1324]), .O(
        n29050) );
  ND2S U31130 ( .I1(n29124), .I2(img[1388]), .O(n29049) );
  ND3S U31131 ( .I1(n29197), .I2(n29050), .I3(n29049), .O(n29052) );
  MUX2 U31132 ( .A(img[1364]), .B(n29052), .S(n29051), .O(n12168) );
  AOI22S U31133 ( .A1(n29072), .A2(img[1388]), .B1(n13781), .B2(n31877), .O(
        n29053) );
  ND2S U31134 ( .I1(n13806), .I2(n29053), .O(n29055) );
  MUX2 U31135 ( .A(n29055), .B(img[1300]), .S(n29054), .O(n12232) );
  AOI22S U31136 ( .A1(n13779), .A2(n31878), .B1(n29257), .B2(img[1300]), .O(
        n29057) );
  ND2S U31137 ( .I1(n29124), .I2(img[1364]), .O(n29056) );
  ND3S U31138 ( .I1(n29197), .I2(n29057), .I3(n29056), .O(n29059) );
  MUX2 U31139 ( .A(img[1388]), .B(n29059), .S(n29058), .O(n12144) );
  AOI22S U31140 ( .A1(n29072), .A2(img[1004]), .B1(n28913), .B2(n31879), .O(
        n29060) );
  ND2S U31141 ( .I1(n13806), .I2(n29060), .O(n29062) );
  AOI22S U31142 ( .A1(n29072), .A2(img[916]), .B1(n29407), .B2(n31880), .O(
        n29063) );
  ND2S U31143 ( .I1(n13806), .I2(n29063), .O(n29065) );
  MUX2 U31144 ( .A(img[1004]), .B(n29065), .S(n29064), .O(n12528) );
  AOI22S U31145 ( .A1(n29072), .A2(img[236]), .B1(n25859), .B2(n31881), .O(
        n29066) );
  ND2S U31146 ( .I1(n13806), .I2(n29066), .O(n29068) );
  MUX2 U31147 ( .A(img[148]), .B(n29068), .S(n29067), .O(n13384) );
  AOI22S U31148 ( .A1(n29072), .A2(img[148]), .B1(n24193), .B2(n31882), .O(
        n29069) );
  ND2S U31149 ( .I1(n13806), .I2(n29069), .O(n29071) );
  MUX2 U31150 ( .A(img[236]), .B(n29071), .S(n29070), .O(n13296) );
  AOI22S U31151 ( .A1(n29072), .A2(img[364]), .B1(n28862), .B2(n31883), .O(
        n29073) );
  ND2S U31152 ( .I1(n13806), .I2(n29073), .O(n29075) );
  AOI22S U31153 ( .A1(n28442), .A2(img[276]), .B1(n29530), .B2(n31884), .O(
        n29077) );
  ND2S U31154 ( .I1(n13806), .I2(n29077), .O(n29079) );
  MUX2 U31155 ( .A(img[364]), .B(n29079), .S(n29078), .O(n13168) );
  AOI22S U31156 ( .A1(n26970), .A2(img[492]), .B1(n23941), .B2(n31885), .O(
        n29080) );
  ND2S U31157 ( .I1(n13806), .I2(n29080), .O(n29082) );
  AOI22S U31158 ( .A1(n13771), .A2(img[404]), .B1(n28075), .B2(n31886), .O(
        n29083) );
  ND2S U31159 ( .I1(n13806), .I2(n29083), .O(n29085) );
  MUX2 U31160 ( .A(img[492]), .B(n29085), .S(n29084), .O(n13040) );
  AOI22S U31161 ( .A1(n26855), .A2(img[1492]), .B1(n28343), .B2(n31887), .O(
        n29086) );
  ND2S U31162 ( .I1(n13806), .I2(n29086), .O(n29088) );
  AOI22S U31163 ( .A1(n29096), .A2(n31888), .B1(n24313), .B2(img[1452]), .O(
        n29090) );
  ND2S U31164 ( .I1(n29124), .I2(img[1516]), .O(n29089) );
  ND3S U31165 ( .I1(n29197), .I2(n29090), .I3(n29089), .O(n29092) );
  MUX2 U31166 ( .A(n29092), .B(img[1492]), .S(n29091), .O(n12040) );
  AOI22S U31167 ( .A1(n28318), .A2(img[1516]), .B1(n28862), .B2(n31889), .O(
        n29093) );
  ND2S U31168 ( .I1(n13806), .I2(n29093), .O(n29095) );
  MUX2 U31169 ( .A(img[1428]), .B(n29095), .S(n29094), .O(n12104) );
  AOI22S U31170 ( .A1(n29096), .A2(n31890), .B1(n28069), .B2(img[1428]), .O(
        n29098) );
  ND3S U31171 ( .I1(n29197), .I2(n29098), .I3(n29097), .O(n29100) );
  AOI22S U31172 ( .A1(n28318), .A2(img[876]), .B1(n28037), .B2(n31891), .O(
        n29101) );
  ND2S U31173 ( .I1(n13806), .I2(n29101), .O(n29103) );
  INV1S U31174 ( .I(img[876]), .O(n29104) );
  AOI22S U31175 ( .A1(n28318), .A2(img[788]), .B1(n28343), .B2(n29104), .O(
        n29105) );
  ND2S U31176 ( .I1(n13806), .I2(n29105), .O(n29107) );
  AOI22S U31177 ( .A1(n28318), .A2(img[748]), .B1(n28075), .B2(n31892), .O(
        n29108) );
  ND2S U31178 ( .I1(n13806), .I2(n29108), .O(n29110) );
  AOI22S U31179 ( .A1(n28318), .A2(img[660]), .B1(n25062), .B2(n31893), .O(
        n29111) );
  ND2S U31180 ( .I1(n29197), .I2(n29111), .O(n29113) );
  AOI22S U31181 ( .A1(n28318), .A2(img[1108]), .B1(n28862), .B2(n31894), .O(
        n29114) );
  ND2S U31182 ( .I1(n29197), .I2(n29114), .O(n29116) );
  MUX2 U31183 ( .A(n29116), .B(img[1068]), .S(n29115), .O(n12464) );
  AOI22S U31184 ( .A1(n28938), .A2(n31895), .B1(n24313), .B2(img[1068]), .O(
        n29118) );
  ND2S U31185 ( .I1(n29124), .I2(img[1132]), .O(n29117) );
  ND3S U31186 ( .I1(n29197), .I2(n29118), .I3(n29117), .O(n29120) );
  MUX2 U31187 ( .A(img[1108]), .B(n29120), .S(n29119), .O(n12424) );
  AOI22S U31188 ( .A1(n28318), .A2(img[1132]), .B1(n27735), .B2(n31896), .O(
        n29121) );
  ND2S U31189 ( .I1(n29197), .I2(n29121), .O(n29123) );
  MUX2 U31190 ( .A(n29123), .B(img[1044]), .S(n29122), .O(n12487) );
  AOI22S U31191 ( .A1(n13781), .A2(n31897), .B1(n28254), .B2(img[1044]), .O(
        n29126) );
  ND2S U31192 ( .I1(n29124), .I2(img[1108]), .O(n29125) );
  ND3S U31193 ( .I1(n29197), .I2(n29126), .I3(n29125), .O(n29128) );
  MUX2 U31194 ( .A(img[1132]), .B(n29128), .S(n29127), .O(n12400) );
  AOI22S U31195 ( .A1(n29414), .A2(img[596]), .B1(n28862), .B2(n31898), .O(
        n29130) );
  ND2S U31196 ( .I1(n13806), .I2(n29130), .O(n29131) );
  MUX2 U31197 ( .A(n29131), .B(img[556]), .S(n29439), .O(n12976) );
  AOI22S U31198 ( .A1(n28840), .A2(img[556]), .B1(n29407), .B2(n31899), .O(
        n29132) );
  ND2S U31199 ( .I1(n29197), .I2(n29132), .O(n29134) );
  MUX2 U31200 ( .A(n29134), .B(img[596]), .S(n29133), .O(n12936) );
  AOI22S U31201 ( .A1(n26855), .A2(img[84]), .B1(n29407), .B2(n31900), .O(
        n29135) );
  ND2S U31202 ( .I1(n29197), .I2(n29135), .O(n29137) );
  AOI22S U31203 ( .A1(n28347), .A2(img[44]), .B1(n24755), .B2(n31901), .O(
        n29138) );
  ND2S U31204 ( .I1(n29197), .I2(n29138), .O(n29140) );
  MUX2 U31205 ( .A(img[84]), .B(n29140), .S(n29139), .O(n13448) );
  AOI22S U31206 ( .A1(n26101), .A2(img[980]), .B1(n29407), .B2(n31902), .O(
        n29141) );
  ND2S U31207 ( .I1(n29197), .I2(n29141), .O(n29143) );
  AOI22S U31208 ( .A1(n28442), .A2(img[940]), .B1(n29530), .B2(n31903), .O(
        n29144) );
  ND2S U31209 ( .I1(n29197), .I2(n29144), .O(n29146) );
  MUX2 U31210 ( .A(img[980]), .B(n29146), .S(n29145), .O(n12552) );
  AOI22S U31211 ( .A1(n27990), .A2(img[212]), .B1(n27049), .B2(n31904), .O(
        n29147) );
  ND2S U31212 ( .I1(n29197), .I2(n29147), .O(n29149) );
  MUX2 U31213 ( .A(img[172]), .B(n29149), .S(n29148), .O(n13360) );
  AOI22S U31214 ( .A1(n25810), .A2(img[172]), .B1(n24755), .B2(n31905), .O(
        n29150) );
  ND2S U31215 ( .I1(n29197), .I2(n29150), .O(n29152) );
  MUX2 U31216 ( .A(img[212]), .B(n29152), .S(n29151), .O(n13320) );
  AOI22S U31217 ( .A1(n27065), .A2(img[340]), .B1(n29407), .B2(n31906), .O(
        n29153) );
  ND2S U31218 ( .I1(n29197), .I2(n29153), .O(n29155) );
  MUX2 U31219 ( .A(img[300]), .B(n29155), .S(n29154), .O(n13232) );
  AOI22S U31220 ( .A1(n28347), .A2(img[300]), .B1(n29397), .B2(n31907), .O(
        n29156) );
  ND2S U31221 ( .I1(n29197), .I2(n29156), .O(n29158) );
  AOI22S U31222 ( .A1(n27746), .A2(img[468]), .B1(n13781), .B2(n31908), .O(
        n29159) );
  ND2S U31223 ( .I1(n29197), .I2(n29159), .O(n29161) );
  MUX2 U31224 ( .A(img[428]), .B(n29161), .S(n29160), .O(n13104) );
  AOI22S U31225 ( .A1(n26855), .A2(img[428]), .B1(n27049), .B2(n31909), .O(
        n29162) );
  ND2S U31226 ( .I1(n29197), .I2(n29162), .O(n29164) );
  AOI22S U31227 ( .A1(n13780), .A2(img[852]), .B1(n29397), .B2(n31910), .O(
        n29165) );
  ND2S U31228 ( .I1(n29197), .I2(n29165), .O(n29167) );
  INV1S U31229 ( .I(img[852]), .O(n29168) );
  AOI22S U31230 ( .A1(n27746), .A2(img[812]), .B1(n28592), .B2(n29168), .O(
        n29169) );
  ND2S U31231 ( .I1(n29197), .I2(n29169), .O(n29171) );
  AOI22S U31232 ( .A1(n27746), .A2(img[724]), .B1(n25062), .B2(n31911), .O(
        n29172) );
  ND2S U31233 ( .I1(n13806), .I2(n29172), .O(n29174) );
  AOI22S U31234 ( .A1(n28442), .A2(img[684]), .B1(n25062), .B2(n31912), .O(
        n29175) );
  ND2S U31235 ( .I1(n29197), .I2(n29175), .O(n29177) );
  AOI22S U31236 ( .A1(n26822), .A2(img[356]), .B1(n28592), .B2(n31913), .O(
        n29178) );
  ND2S U31237 ( .I1(n29197), .I2(n29178), .O(n29180) );
  MUX2 U31238 ( .A(img[284]), .B(n29180), .S(n29179), .O(n13248) );
  AOI22S U31239 ( .A1(n28442), .A2(img[284]), .B1(n29194), .B2(n31914), .O(
        n29181) );
  ND2S U31240 ( .I1(n29197), .I2(n29181), .O(n29183) );
  AOI22S U31241 ( .A1(n27990), .A2(img[1116]), .B1(n28433), .B2(n31915), .O(
        n29184) );
  ND2S U31242 ( .I1(n29197), .I2(n29184), .O(n29186) );
  AOI22S U31243 ( .A1(n29194), .A2(n31916), .B1(n24313), .B2(img[1060]), .O(
        n29188) );
  ND2S U31244 ( .I1(n13903), .I2(img[1124]), .O(n29187) );
  ND3S U31245 ( .I1(n29197), .I2(n29188), .I3(n29187), .O(n29190) );
  MUX2 U31246 ( .A(img[1116]), .B(n29190), .S(n29189), .O(n12416) );
  AOI22S U31247 ( .A1(n26855), .A2(img[1124]), .B1(n25591), .B2(n31917), .O(
        n29191) );
  ND2S U31248 ( .I1(n29197), .I2(n29191), .O(n29193) );
  MUX2 U31249 ( .A(img[1052]), .B(n29193), .S(n29192), .O(n12480) );
  AOI22S U31250 ( .A1(n29194), .A2(n31918), .B1(n24313), .B2(img[1052]), .O(
        n29196) );
  ND3S U31251 ( .I1(n29197), .I2(n29196), .I3(n29195), .O(n29199) );
  MUX2 U31252 ( .A(img[1124]), .B(n29199), .S(n29198), .O(n12408) );
  AOI22S U31253 ( .A1(n28347), .A2(img[740]), .B1(n13781), .B2(n31919), .O(
        n29200) );
  ND2S U31254 ( .I1(n13806), .I2(n29200), .O(n29202) );
  MUX2 U31255 ( .A(img[668]), .B(n29202), .S(n29201), .O(n12864) );
  AOI22S U31256 ( .A1(n28347), .A2(img[668]), .B1(n29457), .B2(n31920), .O(
        n29203) );
  ND2S U31257 ( .I1(n29197), .I2(n29203), .O(n29205) );
  AOI22S U31258 ( .A1(n13776), .A2(img[1244]), .B1(n13775), .B2(n31921), .O(
        n29206) );
  ND2S U31259 ( .I1(n29197), .I2(n29206), .O(n29208) );
  AOI22S U31260 ( .A1(n28862), .A2(n31922), .B1(n29257), .B2(img[1188]), .O(
        n29210) );
  ND3S U31261 ( .I1(n29197), .I2(n29210), .I3(n29209), .O(n29212) );
  MUX2 U31262 ( .A(img[1244]), .B(n29212), .S(n29211), .O(n12288) );
  AOI22S U31263 ( .A1(n28347), .A2(img[1252]), .B1(n13775), .B2(n31923), .O(
        n29213) );
  ND2S U31264 ( .I1(n29197), .I2(n29213), .O(n29215) );
  MUX2 U31265 ( .A(img[1180]), .B(n29215), .S(n29214), .O(n12352) );
  AOI22S U31266 ( .A1(n25468), .A2(n31924), .B1(n29257), .B2(img[1180]), .O(
        n29217) );
  ND3S U31267 ( .I1(n29197), .I2(n29217), .I3(n29216), .O(n29219) );
  MUX2 U31268 ( .A(img[1252]), .B(n29219), .S(n29218), .O(n12280) );
  AOI22S U31269 ( .A1(n13771), .A2(img[996]), .B1(n13775), .B2(n31925), .O(
        n29220) );
  ND2S U31270 ( .I1(n29197), .I2(n29220), .O(n29222) );
  MUX2 U31271 ( .A(img[924]), .B(n29222), .S(n29221), .O(n12608) );
  AOI22S U31272 ( .A1(n29435), .A2(img[924]), .B1(n13775), .B2(n31926), .O(
        n29223) );
  ND2S U31273 ( .I1(n29197), .I2(n29223), .O(n29225) );
  MUX2 U31274 ( .A(img[996]), .B(n29225), .S(n29224), .O(n12536) );
  AOI22S U31275 ( .A1(n29072), .A2(img[868]), .B1(n13775), .B2(n31927), .O(
        n29226) );
  ND2S U31276 ( .I1(n29197), .I2(n29226), .O(n29228) );
  MUX2 U31277 ( .A(img[796]), .B(n29228), .S(n29227), .O(n12736) );
  AOI22S U31278 ( .A1(n26855), .A2(img[796]), .B1(n13775), .B2(n31928), .O(
        n29229) );
  ND2S U31279 ( .I1(n29197), .I2(n29229), .O(n29231) );
  AOI22S U31280 ( .A1(n28442), .A2(img[1372]), .B1(n13775), .B2(n31929), .O(
        n29232) );
  ND2S U31281 ( .I1(n29197), .I2(n29232), .O(n29234) );
  MUX2 U31282 ( .A(n29234), .B(img[1316]), .S(n29233), .O(n12216) );
  AOI22S U31283 ( .A1(n29242), .A2(n31930), .B1(n29257), .B2(img[1316]), .O(
        n29236) );
  ND3S U31284 ( .I1(n29197), .I2(n29236), .I3(n29235), .O(n29238) );
  MUX2 U31285 ( .A(img[1372]), .B(n29238), .S(n29237), .O(n12160) );
  AOI22S U31286 ( .A1(n28840), .A2(img[1380]), .B1(n13775), .B2(n31931), .O(
        n29239) );
  ND2S U31287 ( .I1(n29197), .I2(n29239), .O(n29241) );
  MUX2 U31288 ( .A(img[1308]), .B(n29241), .S(n29240), .O(n12224) );
  AOI22S U31289 ( .A1(n29242), .A2(n31932), .B1(n29257), .B2(img[1308]), .O(
        n29244) );
  ND2S U31290 ( .I1(n29124), .I2(img[1372]), .O(n29243) );
  ND3S U31291 ( .I1(n29197), .I2(n29244), .I3(n29243), .O(n29246) );
  MUX2 U31292 ( .A(img[1380]), .B(n29246), .S(n29245), .O(n12152) );
  AOI22S U31293 ( .A1(n29414), .A2(img[1500]), .B1(n13775), .B2(n31933), .O(
        n29247) );
  ND2S U31294 ( .I1(n29197), .I2(n29247), .O(n29249) );
  MUX2 U31295 ( .A(n29249), .B(img[1444]), .S(n29248), .O(n12088) );
  AOI22S U31296 ( .A1(n27049), .A2(n31934), .B1(n29257), .B2(img[1444]), .O(
        n29251) );
  ND3S U31297 ( .I1(n29197), .I2(n29251), .I3(n29250), .O(n29253) );
  AOI22S U31298 ( .A1(n27990), .A2(img[1508]), .B1(n13775), .B2(n31935), .O(
        n29254) );
  ND2S U31299 ( .I1(n29197), .I2(n29254), .O(n29256) );
  MUX2 U31300 ( .A(n29256), .B(img[1436]), .S(n29255), .O(n12096) );
  AOI22S U31301 ( .A1(n13781), .A2(n31936), .B1(n29257), .B2(img[1436]), .O(
        n29260) );
  ND3S U31302 ( .I1(n29197), .I2(n29260), .I3(n29259), .O(n29262) );
  MUX2 U31303 ( .A(img[1508]), .B(n29262), .S(n29261), .O(n12024) );
  AOI22S U31304 ( .A1(n26822), .A2(img[228]), .B1(n13775), .B2(n31937), .O(
        n29263) );
  ND2S U31305 ( .I1(n29197), .I2(n29263), .O(n29265) );
  MUX2 U31306 ( .A(img[156]), .B(n29265), .S(n29264), .O(n13376) );
  AOI22S U31307 ( .A1(n28382), .A2(img[156]), .B1(n28433), .B2(n31938), .O(
        n29266) );
  ND2S U31308 ( .I1(n13806), .I2(n29266), .O(n29268) );
  MUX2 U31309 ( .A(img[228]), .B(n29268), .S(n29267), .O(n13304) );
  AOI22S U31310 ( .A1(n27990), .A2(img[484]), .B1(n13781), .B2(n31939), .O(
        n29269) );
  ND2S U31311 ( .I1(n29197), .I2(n29269), .O(n29271) );
  MUX2 U31312 ( .A(img[412]), .B(n29271), .S(n29270), .O(n13120) );
  AOI22S U31313 ( .A1(n27990), .A2(img[412]), .B1(n13781), .B2(n31940), .O(
        n29272) );
  ND2S U31314 ( .I1(n29197), .I2(n29272), .O(n29274) );
  AOI22S U31315 ( .A1(n29414), .A2(img[100]), .B1(n13781), .B2(n31941), .O(
        n29275) );
  ND2S U31316 ( .I1(n29197), .I2(n29275), .O(n29277) );
  MUX2 U31317 ( .A(img[28]), .B(n29277), .S(n29276), .O(n13504) );
  BUF2 U31318 ( .I(n29278), .O(n29354) );
  AOI22S U31319 ( .A1(n29072), .A2(img[28]), .B1(n13781), .B2(n31942), .O(
        n29279) );
  ND2S U31320 ( .I1(n29354), .I2(n29279), .O(n29281) );
  MUX2 U31321 ( .A(img[100]), .B(n29281), .S(n29280), .O(n13432) );
  AOI22S U31322 ( .A1(n29072), .A2(img[612]), .B1(n13781), .B2(n31943), .O(
        n29282) );
  ND2S U31323 ( .I1(n29354), .I2(n29282), .O(n29284) );
  MUX2 U31324 ( .A(img[540]), .B(n29284), .S(n29283), .O(n12992) );
  AOI22S U31325 ( .A1(n28382), .A2(img[540]), .B1(n13781), .B2(n31944), .O(
        n29285) );
  ND2S U31326 ( .I1(n29354), .I2(n29285), .O(n29287) );
  MUX2 U31327 ( .A(n29287), .B(img[612]), .S(n29286), .O(n12920) );
  AOI22S U31328 ( .A1(n13771), .A2(img[628]), .B1(n13781), .B2(n31945), .O(
        n29288) );
  ND2S U31329 ( .I1(n29354), .I2(n29288), .O(n29290) );
  AOI22S U31330 ( .A1(n28442), .A2(img[524]), .B1(n13781), .B2(n31946), .O(
        n29291) );
  ND2S U31331 ( .I1(n29354), .I2(n29291), .O(n29293) );
  MUX2 U31332 ( .A(n29293), .B(img[628]), .S(n29292), .O(n12904) );
  AOI22S U31333 ( .A1(n13772), .A2(img[116]), .B1(n13781), .B2(n31947), .O(
        n29294) );
  ND2S U31334 ( .I1(n29354), .I2(n29294), .O(n29296) );
  AOI22S U31335 ( .A1(n13771), .A2(img[12]), .B1(n13781), .B2(n31948), .O(
        n29297) );
  ND2S U31336 ( .I1(n29354), .I2(n29297), .O(n29298) );
  MUX2 U31337 ( .A(img[116]), .B(n29298), .S(n29536), .O(n13416) );
  AOI22S U31338 ( .A1(n28382), .A2(img[1012]), .B1(n13781), .B2(n31949), .O(
        n29299) );
  ND2S U31339 ( .I1(n29354), .I2(n29299), .O(n29301) );
  AOI22S U31340 ( .A1(n27110), .A2(img[908]), .B1(n13781), .B2(n31950), .O(
        n29302) );
  ND2S U31341 ( .I1(n29354), .I2(n29302), .O(n29304) );
  MUX2 U31342 ( .A(img[1012]), .B(n29304), .S(n29303), .O(n12520) );
  AOI22S U31343 ( .A1(n27957), .A2(img[244]), .B1(n29397), .B2(n31951), .O(
        n29305) );
  ND2S U31344 ( .I1(n29354), .I2(n29305), .O(n29307) );
  AOI22S U31345 ( .A1(n28318), .A2(img[140]), .B1(n27049), .B2(n31952), .O(
        n29308) );
  ND2S U31346 ( .I1(n29354), .I2(n29308), .O(n29310) );
  MUX2 U31347 ( .A(img[244]), .B(n29310), .S(n29309), .O(n13288) );
  AOI22S U31348 ( .A1(n28083), .A2(img[372]), .B1(n28862), .B2(n31953), .O(
        n29311) );
  ND2S U31349 ( .I1(n29354), .I2(n29311), .O(n29313) );
  MUX2 U31350 ( .A(n29313), .B(img[268]), .S(n29312), .O(n13264) );
  AOI22S U31351 ( .A1(n27746), .A2(img[268]), .B1(n28862), .B2(n31954), .O(
        n29314) );
  ND2S U31352 ( .I1(n29354), .I2(n29314), .O(n29316) );
  AOI22S U31353 ( .A1(n13773), .A2(img[500]), .B1(n24755), .B2(n31955), .O(
        n29317) );
  ND2S U31354 ( .I1(n29354), .I2(n29317), .O(n29319) );
  MUX2 U31355 ( .A(n29319), .B(img[396]), .S(n29318), .O(n13136) );
  AOI22S U31356 ( .A1(n27746), .A2(img[396]), .B1(n13781), .B2(n31956), .O(
        n29320) );
  ND2S U31357 ( .I1(n29354), .I2(n29320), .O(n29322) );
  MUX2 U31358 ( .A(img[500]), .B(n29322), .S(n29321), .O(n13032) );
  AOI22S U31359 ( .A1(n29414), .A2(img[884]), .B1(n13781), .B2(n31957), .O(
        n29323) );
  ND2S U31360 ( .I1(n29354), .I2(n29323), .O(n29325) );
  INV1S U31361 ( .I(img[884]), .O(n29326) );
  AOI22S U31362 ( .A1(n27746), .A2(img[780]), .B1(n29457), .B2(n29326), .O(
        n29327) );
  ND2S U31363 ( .I1(n29354), .I2(n29327), .O(n29329) );
  MUX2 U31364 ( .A(n29329), .B(img[884]), .S(n29328), .O(n12648) );
  AOI22S U31365 ( .A1(n28083), .A2(img[756]), .B1(n29194), .B2(n31958), .O(
        n29330) );
  ND2S U31366 ( .I1(n29354), .I2(n29330), .O(n29332) );
  AOI22S U31367 ( .A1(n28442), .A2(img[652]), .B1(n28135), .B2(n31959), .O(
        n29333) );
  ND2S U31368 ( .I1(n29354), .I2(n29333), .O(n29335) );
  AOI22S U31369 ( .A1(n29414), .A2(img[604]), .B1(n24755), .B2(n31960), .O(
        n29336) );
  ND2S U31370 ( .I1(n29354), .I2(n29336), .O(n29337) );
  AOI22S U31371 ( .A1(n26855), .A2(img[36]), .B1(n24755), .B2(n31961), .O(
        n29338) );
  ND2S U31372 ( .I1(n29354), .I2(n29338), .O(n29340) );
  MUX2 U31373 ( .A(img[92]), .B(n29340), .S(n29339), .O(n13440) );
  AOI22S U31374 ( .A1(n29414), .A2(img[92]), .B1(n24755), .B2(n31962), .O(
        n29341) );
  ND2S U31375 ( .I1(n29354), .I2(n29341), .O(n29343) );
  MUX2 U31376 ( .A(img[36]), .B(n29343), .S(n29342), .O(n13496) );
  AOI22S U31377 ( .A1(n28840), .A2(img[932]), .B1(n24755), .B2(n31963), .O(
        n29344) );
  ND2S U31378 ( .I1(n29354), .I2(n29344), .O(n29346) );
  MUX2 U31379 ( .A(img[988]), .B(n29346), .S(n29345), .O(n12544) );
  AOI22S U31380 ( .A1(n28382), .A2(img[988]), .B1(n24755), .B2(n31964), .O(
        n29347) );
  ND2S U31381 ( .I1(n29354), .I2(n29347), .O(n29349) );
  AOI22S U31382 ( .A1(n28347), .A2(img[164]), .B1(n24755), .B2(n31965), .O(
        n29350) );
  ND2S U31383 ( .I1(n29354), .I2(n29350), .O(n29352) );
  MUX2 U31384 ( .A(img[220]), .B(n29352), .S(n29351), .O(n13312) );
  AOI22S U31385 ( .A1(n13771), .A2(img[220]), .B1(n24755), .B2(n31966), .O(
        n29353) );
  ND2S U31386 ( .I1(n29354), .I2(n29353), .O(n29356) );
  MUX2 U31387 ( .A(img[164]), .B(n29356), .S(n29355), .O(n13368) );
  AOI22S U31388 ( .A1(n28318), .A2(img[292]), .B1(n24755), .B2(n31967), .O(
        n29357) );
  ND2S U31389 ( .I1(n29197), .I2(n29357), .O(n29359) );
  MUX2 U31390 ( .A(img[348]), .B(n29359), .S(n29358), .O(n13184) );
  AOI22S U31391 ( .A1(n13773), .A2(img[348]), .B1(n24755), .B2(n31968), .O(
        n29360) );
  ND2S U31392 ( .I1(n29197), .I2(n29360), .O(n29362) );
  AOI22S U31393 ( .A1(n28083), .A2(img[420]), .B1(n28343), .B2(n31969), .O(
        n29363) );
  ND2S U31394 ( .I1(n29197), .I2(n29363), .O(n29365) );
  AOI22S U31395 ( .A1(n13776), .A2(img[476]), .B1(n13781), .B2(n31970), .O(
        n29366) );
  ND2S U31396 ( .I1(n29197), .I2(n29366), .O(n29368) );
  MUX2 U31397 ( .A(img[420]), .B(n29368), .S(n29367), .O(n13112) );
  INV1S U31398 ( .I(img[860]), .O(n29369) );
  AOI22S U31399 ( .A1(n13776), .A2(img[804]), .B1(n25062), .B2(n29369), .O(
        n29370) );
  ND2S U31400 ( .I1(n29197), .I2(n29370), .O(n29372) );
  AOI22S U31401 ( .A1(n13776), .A2(img[860]), .B1(n29397), .B2(n31971), .O(
        n29373) );
  ND2S U31402 ( .I1(n29197), .I2(n29373), .O(n29375) );
  AOI22S U31403 ( .A1(n13776), .A2(img[676]), .B1(n29397), .B2(n31972), .O(
        n29376) );
  ND2S U31404 ( .I1(n29197), .I2(n29376), .O(n29378) );
  AOI22S U31405 ( .A1(n13776), .A2(img[732]), .B1(n29397), .B2(n31973), .O(
        n29379) );
  ND2S U31406 ( .I1(n29197), .I2(n29379), .O(n29381) );
  AOI22S U31407 ( .A1(n13776), .A2(img[636]), .B1(n29397), .B2(n31974), .O(
        n29382) );
  ND2S U31408 ( .I1(n29197), .I2(n29382), .O(n29384) );
  MUX2 U31409 ( .A(n29384), .B(img[516]), .S(n29383), .O(n13016) );
  AOI22S U31410 ( .A1(n13776), .A2(img[516]), .B1(n29397), .B2(n31975), .O(
        n29385) );
  ND2S U31411 ( .I1(n29197), .I2(n29385), .O(n29387) );
  MUX2 U31412 ( .A(n29387), .B(img[636]), .S(n29386), .O(n12896) );
  AOI22S U31413 ( .A1(n13776), .A2(img[124]), .B1(n29397), .B2(n31976), .O(
        n29388) );
  ND2S U31414 ( .I1(n29197), .I2(n29388), .O(n29390) );
  AOI22S U31415 ( .A1(n13776), .A2(img[4]), .B1(n29397), .B2(n31977), .O(
        n29391) );
  ND2S U31416 ( .I1(n29197), .I2(n29391), .O(n29393) );
  MUX2 U31417 ( .A(img[124]), .B(n29393), .S(n29392), .O(n13408) );
  AOI22S U31418 ( .A1(n13776), .A2(img[1020]), .B1(n29397), .B2(n31978), .O(
        n29394) );
  ND2S U31419 ( .I1(n29197), .I2(n29394), .O(n29396) );
  AOI22S U31420 ( .A1(n13776), .A2(img[900]), .B1(n29397), .B2(n31979), .O(
        n29398) );
  ND2S U31421 ( .I1(n29197), .I2(n29398), .O(n29400) );
  AOI22S U31422 ( .A1(n27065), .A2(img[252]), .B1(n29407), .B2(n31980), .O(
        n29401) );
  ND2S U31423 ( .I1(n29197), .I2(n29401), .O(n29403) );
  MUX2 U31424 ( .A(n29403), .B(img[132]), .S(n29402), .O(n13400) );
  AOI22S U31425 ( .A1(n29076), .A2(img[132]), .B1(n29407), .B2(n31981), .O(
        n29404) );
  ND2S U31426 ( .I1(n29197), .I2(n29404), .O(n29406) );
  MUX2 U31427 ( .A(img[252]), .B(n29406), .S(n29405), .O(n13279) );
  AOI22S U31428 ( .A1(n28840), .A2(img[380]), .B1(n29407), .B2(n31982), .O(
        n29408) );
  ND2S U31429 ( .I1(n29197), .I2(n29408), .O(n29410) );
  AOI22S U31430 ( .A1(n29435), .A2(img[260]), .B1(n29457), .B2(n31983), .O(
        n29411) );
  ND2S U31431 ( .I1(n29197), .I2(n29411), .O(n29413) );
  MUX2 U31432 ( .A(img[380]), .B(n29413), .S(n29412), .O(n13152) );
  AOI22S U31433 ( .A1(n29435), .A2(img[508]), .B1(n29457), .B2(n31984), .O(
        n29415) );
  ND2S U31434 ( .I1(n29197), .I2(n29415), .O(n29417) );
  INV1S U31435 ( .I(img[508]), .O(n29418) );
  AOI22S U31436 ( .A1(n29435), .A2(img[388]), .B1(n29457), .B2(n29418), .O(
        n29419) );
  ND2S U31437 ( .I1(n29197), .I2(n29419), .O(n29421) );
  MUX2 U31438 ( .A(n29421), .B(img[508]), .S(n29420), .O(n13024) );
  AOI22S U31439 ( .A1(n29435), .A2(img[892]), .B1(n29457), .B2(n31985), .O(
        n29422) );
  ND2S U31440 ( .I1(n29197), .I2(n29422), .O(n29424) );
  INV1S U31441 ( .I(img[892]), .O(n29425) );
  AOI22S U31442 ( .A1(n29435), .A2(img[772]), .B1(n29457), .B2(n29425), .O(
        n29426) );
  ND2S U31443 ( .I1(n29197), .I2(n29426), .O(n29428) );
  AOI22S U31444 ( .A1(n29435), .A2(img[764]), .B1(n29457), .B2(n31986), .O(
        n29429) );
  ND2S U31445 ( .I1(n29197), .I2(n29429), .O(n29431) );
  AOI22S U31446 ( .A1(n29435), .A2(img[644]), .B1(n29457), .B2(n31987), .O(
        n29432) );
  ND2S U31447 ( .I1(n29197), .I2(n29432), .O(n29434) );
  INV1S U31448 ( .I(n29526), .O(n29534) );
  MUX2S U31449 ( .A(A67_shift[12]), .B(A67_shift[4]), .S(n29534), .O(n11388)
         );
  MUX2S U31450 ( .A(A67_shift[20]), .B(A67_shift[12]), .S(n13774), .O(n11387)
         );
  MUX2S U31451 ( .A(A67_shift[28]), .B(A67_shift[20]), .S(n13821), .O(n11386)
         );
  MUX2S U31452 ( .A(A67_shift[36]), .B(A67_shift[28]), .S(n13774), .O(n11385)
         );
  MUX2S U31453 ( .A(A67_shift[44]), .B(A67_shift[36]), .S(n13821), .O(n11384)
         );
  MUX2S U31454 ( .A(A67_shift[52]), .B(A67_shift[44]), .S(n13774), .O(n11383)
         );
  MUX2S U31455 ( .A(A67_shift[60]), .B(A67_shift[52]), .S(n13821), .O(n11382)
         );
  MUX2S U31456 ( .A(A67_shift[68]), .B(A67_shift[60]), .S(n13774), .O(n11381)
         );
  MUX2S U31457 ( .A(A67_shift[76]), .B(A67_shift[68]), .S(n13821), .O(n11380)
         );
  MUX2S U31458 ( .A(A67_shift[84]), .B(A67_shift[76]), .S(n13774), .O(n11379)
         );
  MUX2S U31459 ( .A(A67_shift[92]), .B(A67_shift[84]), .S(n13821), .O(n11378)
         );
  MUX2S U31460 ( .A(A67_shift[100]), .B(A67_shift[92]), .S(n13821), .O(n11377)
         );
  MUX2S U31461 ( .A(A67_shift[108]), .B(A67_shift[100]), .S(n13821), .O(n11376) );
  MUX2S U31462 ( .A(A67_shift[116]), .B(A67_shift[108]), .S(n13821), .O(n11375) );
  MUX2S U31463 ( .A(A67_shift[124]), .B(A67_shift[116]), .S(n13821), .O(n11374) );
  MUX2S U31464 ( .A(A67_shift[132]), .B(A67_shift[124]), .S(n13821), .O(n11373) );
  MUX2S U31465 ( .A(A67_shift[140]), .B(A67_shift[132]), .S(n13821), .O(n11372) );
  MUX2S U31466 ( .A(A67_shift[148]), .B(A67_shift[140]), .S(n13821), .O(n11371) );
  MUX2S U31467 ( .A(A67_shift[156]), .B(A67_shift[148]), .S(n13821), .O(n11370) );
  MUX2S U31468 ( .A(A67_shift[164]), .B(A67_shift[156]), .S(n13821), .O(n11369) );
  MUX2S U31469 ( .A(A67_shift[172]), .B(A67_shift[164]), .S(n13821), .O(n11368) );
  MUX2S U31470 ( .A(A67_shift[180]), .B(A67_shift[172]), .S(n13821), .O(n11367) );
  MUX2S U31471 ( .A(A67_shift[188]), .B(A67_shift[180]), .S(n13821), .O(n11366) );
  MUX2S U31472 ( .A(A67_shift[196]), .B(A67_shift[188]), .S(n13821), .O(n11365) );
  MUX2S U31473 ( .A(A67_shift[204]), .B(A67_shift[196]), .S(n13821), .O(n11364) );
  MUX2S U31474 ( .A(A67_shift[212]), .B(A67_shift[204]), .S(n13821), .O(n11363) );
  MUX2S U31475 ( .A(A67_shift[220]), .B(A67_shift[212]), .S(n13821), .O(n11362) );
  MUX2S U31476 ( .A(A67_shift[228]), .B(A67_shift[220]), .S(n13821), .O(n11361) );
  MUX2S U31477 ( .A(A67_shift[236]), .B(A67_shift[228]), .S(n13821), .O(n11360) );
  MUX2S U31478 ( .A(A67_shift[244]), .B(A67_shift[236]), .S(n13821), .O(n11359) );
  MUX2S U31479 ( .A(A67_shift[252]), .B(A67_shift[244]), .S(n13821), .O(n11358) );
  AOI22S U31480 ( .A1(n29435), .A2(img[548]), .B1(n29457), .B2(n31988), .O(
        n29436) );
  ND2S U31481 ( .I1(n29197), .I2(n29436), .O(n29437) );
  MUX2 U31482 ( .A(n29437), .B(img[604]), .S(n29478), .O(n12928) );
  MUX2S U31483 ( .A(A67_shift[8]), .B(A67_shift[0]), .S(n13821), .O(n11260) );
  MUX2S U31484 ( .A(A67_shift[16]), .B(A67_shift[8]), .S(n13774), .O(n11259)
         );
  MUX2S U31485 ( .A(A67_shift[24]), .B(A67_shift[16]), .S(n13821), .O(n11258)
         );
  MUX2S U31486 ( .A(A67_shift[32]), .B(A67_shift[24]), .S(n13821), .O(n11257)
         );
  MUX2S U31487 ( .A(A67_shift[40]), .B(A67_shift[32]), .S(n13821), .O(n11256)
         );
  MUX2S U31488 ( .A(A67_shift[48]), .B(A67_shift[40]), .S(n13821), .O(n11255)
         );
  MUX2S U31489 ( .A(A67_shift[56]), .B(A67_shift[48]), .S(n13821), .O(n11254)
         );
  MUX2S U31490 ( .A(A67_shift[64]), .B(A67_shift[56]), .S(n13774), .O(n11253)
         );
  MUX2S U31491 ( .A(A67_shift[72]), .B(A67_shift[64]), .S(n13821), .O(n11252)
         );
  MUX2S U31492 ( .A(A67_shift[80]), .B(A67_shift[72]), .S(n13821), .O(n11251)
         );
  MUX2S U31493 ( .A(A67_shift[88]), .B(A67_shift[80]), .S(n13821), .O(n11250)
         );
  MUX2S U31494 ( .A(A67_shift[96]), .B(A67_shift[88]), .S(n13821), .O(n11249)
         );
  MUX2S U31495 ( .A(A67_shift[104]), .B(A67_shift[96]), .S(n13821), .O(n11248)
         );
  MUX2S U31496 ( .A(A67_shift[112]), .B(A67_shift[104]), .S(n13774), .O(n11247) );
  MUX2S U31497 ( .A(A67_shift[120]), .B(A67_shift[112]), .S(n13821), .O(n11246) );
  MUX2S U31498 ( .A(A67_shift[128]), .B(A67_shift[120]), .S(n13821), .O(n11245) );
  MUX2S U31499 ( .A(A67_shift[136]), .B(A67_shift[128]), .S(n13821), .O(n11244) );
  MUX2S U31500 ( .A(A67_shift[144]), .B(A67_shift[136]), .S(n13821), .O(n11243) );
  MUX2S U31501 ( .A(A67_shift[152]), .B(A67_shift[144]), .S(n13821), .O(n11242) );
  MUX2S U31502 ( .A(A67_shift[160]), .B(A67_shift[152]), .S(n13774), .O(n11241) );
  MUX2S U31503 ( .A(A67_shift[168]), .B(A67_shift[160]), .S(n13821), .O(n11240) );
  MUX2S U31504 ( .A(A67_shift[176]), .B(A67_shift[168]), .S(n13774), .O(n11239) );
  MUX2S U31505 ( .A(A67_shift[184]), .B(A67_shift[176]), .S(n13821), .O(n11238) );
  MUX2S U31506 ( .A(A67_shift[192]), .B(A67_shift[184]), .S(n13774), .O(n11237) );
  MUX2S U31507 ( .A(A67_shift[200]), .B(A67_shift[192]), .S(n13821), .O(n11236) );
  MUX2S U31508 ( .A(A67_shift[208]), .B(A67_shift[200]), .S(n13774), .O(n11235) );
  MUX2S U31509 ( .A(A67_shift[216]), .B(A67_shift[208]), .S(n13821), .O(n11234) );
  MUX2S U31510 ( .A(A67_shift[224]), .B(A67_shift[216]), .S(n13774), .O(n11233) );
  MUX2S U31511 ( .A(A67_shift[232]), .B(A67_shift[224]), .S(n13821), .O(n11232) );
  MUX2S U31512 ( .A(A67_shift[240]), .B(A67_shift[232]), .S(n13774), .O(n11231) );
  MUX2S U31513 ( .A(A67_shift[248]), .B(A67_shift[240]), .S(n13821), .O(n11229) );
  AOI22S U31514 ( .A1(n27746), .A2(img[592]), .B1(n29457), .B2(n31989), .O(
        n29438) );
  ND2S U31515 ( .I1(n28425), .I2(n29438), .O(n29440) );
  MUX2 U31516 ( .A(n29440), .B(img[552]), .S(n29439), .O(n12980) );
  MOAI1 U31517 ( .A1(n29504), .A2(n29442), .B1(n29502), .B2(n29441), .O(n29454) );
  AOI22S U31518 ( .A1(n29507), .A2(n29444), .B1(n29506), .B2(n29443), .O(
        n29447) );
  ND2S U31519 ( .I1(n29510), .I2(n29445), .O(n29446) );
  OAI112HS U31520 ( .C1(n29514), .C2(n29448), .A1(n29447), .B1(n29446), .O(
        n29449) );
  AOI13HS U31521 ( .B1(n29518), .B2(n29450), .B3(n29516), .A1(n29449), .O(
        n29453) );
  ND2 U31522 ( .I1(n29521), .I2(n29451), .O(n29452) );
  OR3B2 U31523 ( .I1(n29454), .B1(n29453), .B2(n29452), .O(n29456) );
  AO222 U31524 ( .A1(n29456), .A2(n29527), .B1(n29526), .B2(A67_shift[3]), 
        .C1(n29455), .C2(n29525), .O(n11357) );
  MUX2S U31525 ( .A(A67_shift[11]), .B(A67_shift[3]), .S(n13774), .O(n11356)
         );
  MUX2S U31526 ( .A(A67_shift[19]), .B(A67_shift[11]), .S(n13821), .O(n11355)
         );
  MUX2S U31527 ( .A(A67_shift[27]), .B(A67_shift[19]), .S(n29529), .O(n11354)
         );
  MUX2S U31528 ( .A(A67_shift[35]), .B(A67_shift[27]), .S(n29529), .O(n11353)
         );
  MUX2S U31529 ( .A(A67_shift[43]), .B(A67_shift[35]), .S(n29534), .O(n11352)
         );
  MUX2S U31530 ( .A(A67_shift[51]), .B(A67_shift[43]), .S(n29529), .O(n11351)
         );
  MUX2S U31531 ( .A(A67_shift[59]), .B(A67_shift[51]), .S(n29534), .O(n11350)
         );
  MUX2S U31532 ( .A(A67_shift[67]), .B(A67_shift[59]), .S(n29529), .O(n11349)
         );
  MUX2S U31533 ( .A(A67_shift[75]), .B(A67_shift[67]), .S(n13774), .O(n11348)
         );
  MUX2S U31534 ( .A(A67_shift[83]), .B(A67_shift[75]), .S(n13774), .O(n11347)
         );
  MUX2S U31535 ( .A(A67_shift[91]), .B(A67_shift[83]), .S(n13774), .O(n11346)
         );
  MUX2S U31536 ( .A(A67_shift[99]), .B(A67_shift[91]), .S(n13774), .O(n11345)
         );
  MUX2S U31537 ( .A(A67_shift[107]), .B(A67_shift[99]), .S(n13774), .O(n11344)
         );
  MUX2S U31538 ( .A(A67_shift[115]), .B(A67_shift[107]), .S(n13774), .O(n11343) );
  MUX2S U31539 ( .A(A67_shift[123]), .B(A67_shift[115]), .S(n13774), .O(n11342) );
  MUX2S U31540 ( .A(A67_shift[131]), .B(A67_shift[123]), .S(n13774), .O(n11341) );
  MUX2S U31541 ( .A(A67_shift[139]), .B(A67_shift[131]), .S(n13774), .O(n11340) );
  MUX2S U31542 ( .A(A67_shift[147]), .B(A67_shift[139]), .S(n13774), .O(n11339) );
  MUX2S U31543 ( .A(A67_shift[155]), .B(A67_shift[147]), .S(n13774), .O(n11338) );
  MUX2S U31544 ( .A(A67_shift[163]), .B(A67_shift[155]), .S(n13774), .O(n11337) );
  MUX2S U31545 ( .A(A67_shift[171]), .B(A67_shift[163]), .S(n13774), .O(n11336) );
  MUX2S U31546 ( .A(A67_shift[179]), .B(A67_shift[171]), .S(n13774), .O(n11335) );
  MUX2S U31547 ( .A(A67_shift[187]), .B(A67_shift[179]), .S(n13774), .O(n11334) );
  MUX2S U31548 ( .A(A67_shift[195]), .B(A67_shift[187]), .S(n13774), .O(n11333) );
  MUX2S U31549 ( .A(A67_shift[203]), .B(A67_shift[195]), .S(n13774), .O(n11332) );
  MUX2S U31550 ( .A(A67_shift[211]), .B(A67_shift[203]), .S(n13774), .O(n11331) );
  MUX2S U31551 ( .A(A67_shift[219]), .B(A67_shift[211]), .S(n13774), .O(n11330) );
  MUX2S U31552 ( .A(A67_shift[227]), .B(A67_shift[219]), .S(n13774), .O(n11329) );
  MUX2S U31553 ( .A(A67_shift[235]), .B(A67_shift[227]), .S(n13774), .O(n11328) );
  MUX2S U31554 ( .A(A67_shift[243]), .B(A67_shift[235]), .S(n13774), .O(n11327) );
  MUX2S U31555 ( .A(A67_shift[251]), .B(A67_shift[243]), .S(n13821), .O(n11326) );
  AOI22S U31556 ( .A1(n27746), .A2(img[603]), .B1(n29457), .B2(n31990), .O(
        n29458) );
  ND2S U31557 ( .I1(n27886), .I2(n29458), .O(n29459) );
  MOAI1 U31558 ( .A1(n29504), .A2(n29461), .B1(n29502), .B2(n29460), .O(n29474) );
  AOI22S U31559 ( .A1(n29507), .A2(n29463), .B1(n29506), .B2(n29462), .O(
        n29466) );
  OAI112HS U31560 ( .C1(n29514), .C2(n29467), .A1(n29466), .B1(n29465), .O(
        n29468) );
  INV1S U31561 ( .I(n29470), .O(n29471) );
  ND2 U31562 ( .I1(n29521), .I2(n29471), .O(n29472) );
  OR3B2 U31563 ( .I1(n29474), .B1(n29473), .B2(n29472), .O(n29476) );
  AO222 U31564 ( .A1(n29476), .A2(n29527), .B1(n29526), .B2(A67_shift[1]), 
        .C1(n29475), .C2(n29525), .O(n11293) );
  MUX2S U31565 ( .A(A67_shift[9]), .B(A67_shift[1]), .S(n13774), .O(n11292) );
  MUX2S U31566 ( .A(A67_shift[17]), .B(A67_shift[9]), .S(n13821), .O(n11291)
         );
  MUX2S U31567 ( .A(A67_shift[25]), .B(A67_shift[17]), .S(n13774), .O(n11290)
         );
  MUX2S U31568 ( .A(A67_shift[33]), .B(A67_shift[25]), .S(n13774), .O(n11289)
         );
  MUX2S U31569 ( .A(A67_shift[41]), .B(A67_shift[33]), .S(n13821), .O(n11288)
         );
  MUX2S U31570 ( .A(A67_shift[49]), .B(A67_shift[41]), .S(n13821), .O(n11287)
         );
  MUX2S U31571 ( .A(A67_shift[57]), .B(A67_shift[49]), .S(n13821), .O(n11286)
         );
  MUX2S U31572 ( .A(A67_shift[65]), .B(A67_shift[57]), .S(n13821), .O(n11285)
         );
  MUX2S U31573 ( .A(A67_shift[73]), .B(A67_shift[65]), .S(n13774), .O(n11284)
         );
  MUX2S U31574 ( .A(A67_shift[81]), .B(A67_shift[73]), .S(n13821), .O(n11283)
         );
  MUX2S U31575 ( .A(A67_shift[89]), .B(A67_shift[81]), .S(n13774), .O(n11282)
         );
  MUX2S U31576 ( .A(A67_shift[97]), .B(A67_shift[89]), .S(n13821), .O(n11281)
         );
  MUX2S U31577 ( .A(A67_shift[105]), .B(A67_shift[97]), .S(n13774), .O(n11280)
         );
  MUX2S U31578 ( .A(A67_shift[113]), .B(A67_shift[105]), .S(n13774), .O(n11279) );
  MUX2S U31579 ( .A(A67_shift[121]), .B(A67_shift[113]), .S(n13821), .O(n11278) );
  MUX2S U31580 ( .A(A67_shift[129]), .B(A67_shift[121]), .S(n13821), .O(n11277) );
  MUX2S U31581 ( .A(A67_shift[137]), .B(A67_shift[129]), .S(n13821), .O(n11276) );
  MUX2S U31582 ( .A(A67_shift[145]), .B(A67_shift[137]), .S(n13774), .O(n11275) );
  MUX2S U31583 ( .A(A67_shift[153]), .B(A67_shift[145]), .S(n29534), .O(n11274) );
  MUX2S U31584 ( .A(A67_shift[161]), .B(A67_shift[153]), .S(n13821), .O(n11273) );
  MUX2S U31585 ( .A(A67_shift[169]), .B(A67_shift[161]), .S(n13774), .O(n11272) );
  MUX2S U31586 ( .A(A67_shift[177]), .B(A67_shift[169]), .S(n23770), .O(n11271) );
  MUX2S U31587 ( .A(A67_shift[185]), .B(A67_shift[177]), .S(n13774), .O(n11270) );
  MUX2S U31588 ( .A(A67_shift[193]), .B(A67_shift[185]), .S(n13774), .O(n11269) );
  MUX2S U31589 ( .A(A67_shift[201]), .B(A67_shift[193]), .S(n23770), .O(n11268) );
  AOI22S U31590 ( .A1(n27065), .A2(img[545]), .B1(n24755), .B2(n31991), .O(
        n29477) );
  ND2S U31591 ( .I1(n27070), .I2(n29477), .O(n29479) );
  MUX2 U31592 ( .A(n29479), .B(img[601]), .S(n29478), .O(n12931) );
  MUX2S U31593 ( .A(A67_shift[13]), .B(A67_shift[5]), .S(n13821), .O(n11420)
         );
  MUX2S U31594 ( .A(A67_shift[21]), .B(A67_shift[13]), .S(n13774), .O(n11419)
         );
  MUX2S U31595 ( .A(A67_shift[29]), .B(A67_shift[21]), .S(n23770), .O(n11418)
         );
  MUX2S U31596 ( .A(A67_shift[37]), .B(A67_shift[29]), .S(n13774), .O(n11417)
         );
  MUX2S U31597 ( .A(A67_shift[45]), .B(A67_shift[37]), .S(n13774), .O(n11416)
         );
  MUX2S U31598 ( .A(A67_shift[53]), .B(A67_shift[45]), .S(n23770), .O(n11415)
         );
  MUX2S U31599 ( .A(A67_shift[61]), .B(A67_shift[53]), .S(n13774), .O(n11414)
         );
  MUX2S U31600 ( .A(A67_shift[69]), .B(A67_shift[61]), .S(n13774), .O(n11413)
         );
  INV1S U31601 ( .I(n29526), .O(n29529) );
  MUX2S U31602 ( .A(A67_shift[77]), .B(A67_shift[69]), .S(n29529), .O(n11412)
         );
  MUX2S U31603 ( .A(A67_shift[85]), .B(A67_shift[77]), .S(n29534), .O(n11411)
         );
  MUX2S U31604 ( .A(A67_shift[93]), .B(A67_shift[85]), .S(n13774), .O(n11410)
         );
  MUX2S U31605 ( .A(A67_shift[101]), .B(A67_shift[93]), .S(n29529), .O(n11409)
         );
  MUX2S U31606 ( .A(A67_shift[109]), .B(A67_shift[101]), .S(n29534), .O(n11408) );
  MUX2S U31607 ( .A(A67_shift[117]), .B(A67_shift[109]), .S(n13774), .O(n11407) );
  MUX2S U31608 ( .A(A67_shift[125]), .B(A67_shift[117]), .S(n29529), .O(n11406) );
  MUX2S U31609 ( .A(A67_shift[133]), .B(A67_shift[125]), .S(n29534), .O(n11405) );
  MUX2S U31610 ( .A(A67_shift[141]), .B(A67_shift[133]), .S(n13774), .O(n11404) );
  MUX2S U31611 ( .A(A67_shift[149]), .B(A67_shift[141]), .S(n29529), .O(n11403) );
  MUX2S U31612 ( .A(A67_shift[157]), .B(A67_shift[149]), .S(n29534), .O(n11402) );
  MUX2S U31613 ( .A(A67_shift[165]), .B(A67_shift[157]), .S(n13774), .O(n11401) );
  MUX2S U31614 ( .A(A67_shift[173]), .B(A67_shift[165]), .S(n29529), .O(n11400) );
  MUX2S U31615 ( .A(A67_shift[181]), .B(A67_shift[173]), .S(n29529), .O(n11399) );
  MUX2S U31616 ( .A(A67_shift[189]), .B(A67_shift[181]), .S(n29529), .O(n11398) );
  MUX2S U31617 ( .A(A67_shift[197]), .B(A67_shift[189]), .S(n29529), .O(n11397) );
  MUX2S U31618 ( .A(A67_shift[205]), .B(A67_shift[197]), .S(n29529), .O(n11396) );
  MUX2S U31619 ( .A(A67_shift[213]), .B(A67_shift[205]), .S(n29529), .O(n11395) );
  MUX2S U31620 ( .A(A67_shift[221]), .B(A67_shift[213]), .S(n29529), .O(n11394) );
  MUX2S U31621 ( .A(A67_shift[229]), .B(A67_shift[221]), .S(n29529), .O(n11393) );
  MUX2S U31622 ( .A(A67_shift[237]), .B(A67_shift[229]), .S(n29529), .O(n11392) );
  MUX2S U31623 ( .A(A67_shift[245]), .B(A67_shift[237]), .S(n29529), .O(n11391) );
  MUX2S U31624 ( .A(A67_shift[253]), .B(A67_shift[245]), .S(n29529), .O(n11390) );
  AOI22S U31625 ( .A1(n13776), .A2(img[605]), .B1(n13781), .B2(n31992), .O(
        n29480) );
  ND2S U31626 ( .I1(n13767), .I2(n29480), .O(n29482) );
  NR2P U31627 ( .I1(n29483), .I2(n29504), .O(n29496) );
  AOI22S U31628 ( .A1(n29507), .A2(n29485), .B1(n29506), .B2(n29484), .O(
        n29488) );
  ND2S U31629 ( .I1(n29510), .I2(n29486), .O(n29487) );
  OR3B2 U31630 ( .I1(n29496), .B1(n29495), .B2(n29494), .O(n29498) );
  AO222 U31631 ( .A1(n29498), .A2(n29527), .B1(n29526), .B2(A67_shift[2]), 
        .C1(n29497), .C2(n29525), .O(n11325) );
  MUX2S U31632 ( .A(A67_shift[10]), .B(A67_shift[2]), .S(n29529), .O(n11324)
         );
  MUX2S U31633 ( .A(A67_shift[18]), .B(A67_shift[10]), .S(n29529), .O(n11323)
         );
  MUX2S U31634 ( .A(A67_shift[26]), .B(A67_shift[18]), .S(n29529), .O(n11322)
         );
  MUX2S U31635 ( .A(A67_shift[34]), .B(A67_shift[26]), .S(n29529), .O(n11321)
         );
  MUX2S U31636 ( .A(A67_shift[42]), .B(A67_shift[34]), .S(n29529), .O(n11320)
         );
  MUX2S U31637 ( .A(A67_shift[50]), .B(A67_shift[42]), .S(n29529), .O(n11319)
         );
  MUX2S U31638 ( .A(A67_shift[58]), .B(A67_shift[50]), .S(n29529), .O(n11318)
         );
  MUX2S U31639 ( .A(A67_shift[66]), .B(A67_shift[58]), .S(n29529), .O(n11317)
         );
  MUX2S U31640 ( .A(A67_shift[74]), .B(A67_shift[66]), .S(n29529), .O(n11316)
         );
  MUX2S U31641 ( .A(A67_shift[82]), .B(A67_shift[74]), .S(n13774), .O(n11315)
         );
  MUX2S U31642 ( .A(A67_shift[90]), .B(A67_shift[82]), .S(n13774), .O(n11314)
         );
  MUX2S U31643 ( .A(A67_shift[98]), .B(A67_shift[90]), .S(n13774), .O(n11313)
         );
  MUX2S U31644 ( .A(A67_shift[106]), .B(A67_shift[98]), .S(n13774), .O(n11312)
         );
  MUX2S U31645 ( .A(A67_shift[114]), .B(A67_shift[106]), .S(n13774), .O(n11311) );
  MUX2S U31646 ( .A(A67_shift[122]), .B(A67_shift[114]), .S(n13774), .O(n11310) );
  MUX2S U31647 ( .A(A67_shift[130]), .B(A67_shift[122]), .S(n13774), .O(n11309) );
  MUX2S U31648 ( .A(A67_shift[138]), .B(A67_shift[130]), .S(n13774), .O(n11308) );
  MUX2S U31649 ( .A(A67_shift[146]), .B(A67_shift[138]), .S(n13774), .O(n11307) );
  MUX2S U31650 ( .A(A67_shift[154]), .B(A67_shift[146]), .S(n13774), .O(n11306) );
  MUX2S U31651 ( .A(A67_shift[162]), .B(A67_shift[154]), .S(n13774), .O(n11305) );
  MUX2S U31652 ( .A(A67_shift[170]), .B(A67_shift[162]), .S(n13774), .O(n11304) );
  MUX2S U31653 ( .A(A67_shift[178]), .B(A67_shift[170]), .S(n13774), .O(n11303) );
  MUX2S U31654 ( .A(A67_shift[186]), .B(A67_shift[178]), .S(n13774), .O(n11302) );
  MUX2S U31655 ( .A(A67_shift[194]), .B(A67_shift[186]), .S(n13774), .O(n11301) );
  MUX2S U31656 ( .A(A67_shift[202]), .B(A67_shift[194]), .S(n13774), .O(n11300) );
  MUX2S U31657 ( .A(A67_shift[210]), .B(A67_shift[202]), .S(n13774), .O(n11299) );
  MUX2S U31658 ( .A(A67_shift[218]), .B(A67_shift[210]), .S(n13774), .O(n11298) );
  MUX2S U31659 ( .A(A67_shift[226]), .B(A67_shift[218]), .S(n13774), .O(n11297) );
  MUX2S U31660 ( .A(A67_shift[234]), .B(A67_shift[226]), .S(n13774), .O(n11296) );
  MUX2S U31661 ( .A(A67_shift[242]), .B(A67_shift[234]), .S(n29529), .O(n11295) );
  MUX2S U31662 ( .A(A67_shift[250]), .B(A67_shift[242]), .S(n29534), .O(n11294) );
  AOI22S U31663 ( .A1(n28840), .A2(img[578]), .B1(n29530), .B2(n31993), .O(
        n29499) );
  ND2S U31664 ( .I1(n26010), .I2(n29499), .O(n29500) );
  MUX2 U31665 ( .A(n29500), .B(img[570]), .S(n29532), .O(n12962) );
  MOAI1 U31666 ( .A1(n29504), .A2(n29503), .B1(n29502), .B2(n29501), .O(n29524) );
  INV1S U31667 ( .I(n17965), .O(n29517) );
  AOI22S U31668 ( .A1(n29508), .A2(n29507), .B1(n29506), .B2(n29505), .O(
        n29512) );
  ND2S U31669 ( .I1(n29510), .I2(n29509), .O(n29511) );
  OAI112HS U31670 ( .C1(n29514), .C2(n29513), .A1(n29512), .B1(n29511), .O(
        n29515) );
  AOI13HS U31671 ( .B1(n29518), .B2(n29517), .B3(n29516), .A1(n29515), .O(
        n29523) );
  INV1S U31672 ( .I(n29519), .O(n29520) );
  ND2 U31673 ( .I1(n29521), .I2(n29520), .O(n29522) );
  OR3B2 U31674 ( .I1(n29524), .B1(n29523), .B2(n29522), .O(n29528) );
  AO222 U31675 ( .A1(n29528), .A2(n29527), .B1(n29526), .B2(A67_shift[6]), 
        .C1(n21416), .C2(n29525), .O(n11453) );
  MUX2S U31676 ( .A(A67_shift[14]), .B(A67_shift[6]), .S(n13774), .O(n11452)
         );
  MUX2S U31677 ( .A(A67_shift[22]), .B(A67_shift[14]), .S(n29529), .O(n11451)
         );
  MUX2S U31678 ( .A(A67_shift[30]), .B(A67_shift[22]), .S(n29534), .O(n11450)
         );
  MUX2S U31679 ( .A(A67_shift[38]), .B(A67_shift[30]), .S(n13774), .O(n11449)
         );
  MUX2S U31680 ( .A(A67_shift[46]), .B(A67_shift[38]), .S(n29529), .O(n11448)
         );
  MUX2S U31681 ( .A(A67_shift[54]), .B(A67_shift[46]), .S(n29534), .O(n11447)
         );
  MUX2S U31682 ( .A(A67_shift[62]), .B(A67_shift[54]), .S(n29529), .O(n11446)
         );
  MUX2S U31683 ( .A(A67_shift[70]), .B(A67_shift[62]), .S(n29534), .O(n11445)
         );
  MUX2S U31684 ( .A(A67_shift[78]), .B(A67_shift[70]), .S(n13774), .O(n11444)
         );
  MUX2S U31685 ( .A(A67_shift[86]), .B(A67_shift[78]), .S(n29529), .O(n11443)
         );
  MUX2S U31686 ( .A(A67_shift[94]), .B(A67_shift[86]), .S(n29534), .O(n11442)
         );
  MUX2S U31687 ( .A(A67_shift[102]), .B(A67_shift[94]), .S(n13774), .O(n11441)
         );
  MUX2S U31688 ( .A(A67_shift[110]), .B(A67_shift[102]), .S(n29529), .O(n11440) );
  MUX2S U31689 ( .A(A67_shift[118]), .B(A67_shift[110]), .S(n29534), .O(n11439) );
  MUX2S U31690 ( .A(A67_shift[126]), .B(A67_shift[118]), .S(n13774), .O(n11438) );
  MUX2S U31691 ( .A(A67_shift[134]), .B(A67_shift[126]), .S(n29529), .O(n11437) );
  MUX2S U31692 ( .A(A67_shift[142]), .B(A67_shift[134]), .S(n29534), .O(n11436) );
  MUX2S U31693 ( .A(A67_shift[150]), .B(A67_shift[142]), .S(n29534), .O(n11435) );
  MUX2S U31694 ( .A(A67_shift[158]), .B(A67_shift[150]), .S(n29534), .O(n11434) );
  MUX2S U31695 ( .A(A67_shift[166]), .B(A67_shift[158]), .S(n29534), .O(n11433) );
  MUX2S U31696 ( .A(A67_shift[174]), .B(A67_shift[166]), .S(n29534), .O(n11432) );
  MUX2S U31697 ( .A(A67_shift[182]), .B(A67_shift[174]), .S(n29534), .O(n11431) );
  MUX2S U31698 ( .A(A67_shift[190]), .B(A67_shift[182]), .S(n29534), .O(n11430) );
  MUX2S U31699 ( .A(A67_shift[198]), .B(A67_shift[190]), .S(n29534), .O(n11429) );
  MUX2S U31700 ( .A(A67_shift[206]), .B(A67_shift[198]), .S(n29534), .O(n11428) );
  MUX2S U31701 ( .A(A67_shift[214]), .B(A67_shift[206]), .S(n29534), .O(n11427) );
  MUX2S U31702 ( .A(A67_shift[222]), .B(A67_shift[214]), .S(n29534), .O(n11426) );
  MUX2S U31703 ( .A(A67_shift[230]), .B(A67_shift[222]), .S(n29534), .O(n11425) );
  MUX2S U31704 ( .A(A67_shift[238]), .B(A67_shift[230]), .S(n29534), .O(n11424) );
  MUX2S U31705 ( .A(A67_shift[246]), .B(A67_shift[238]), .S(n29534), .O(n11423) );
  MUX2S U31706 ( .A(A67_shift[254]), .B(A67_shift[246]), .S(n29534), .O(n11422) );
  AOI22S U31707 ( .A1(n24415), .A2(img[582]), .B1(n29530), .B2(n31994), .O(
        n29531) );
  ND2S U31708 ( .I1(n25327), .I2(n29531), .O(n29533) );
  MUX2 U31709 ( .A(n29533), .B(img[574]), .S(n29532), .O(n12958) );
  MUX2S U31710 ( .A(A67_shift[15]), .B(A67_shift[7]), .S(n29534), .O(n11484)
         );
  MUX2S U31711 ( .A(A67_shift[23]), .B(A67_shift[15]), .S(n29534), .O(n11483)
         );
  MUX2S U31712 ( .A(A67_shift[31]), .B(A67_shift[23]), .S(n29534), .O(n11482)
         );
  MUX2S U31713 ( .A(A67_shift[39]), .B(A67_shift[31]), .S(n29534), .O(n11481)
         );
  MUX2S U31714 ( .A(A67_shift[47]), .B(A67_shift[39]), .S(n29534), .O(n11480)
         );
  MUX2S U31715 ( .A(A67_shift[55]), .B(A67_shift[47]), .S(n29534), .O(n11479)
         );
  MUX2S U31716 ( .A(A67_shift[63]), .B(A67_shift[55]), .S(n13821), .O(n11478)
         );
  MUX2S U31717 ( .A(A67_shift[71]), .B(A67_shift[63]), .S(n13821), .O(n11477)
         );
  MUX2S U31718 ( .A(A67_shift[79]), .B(A67_shift[71]), .S(n13821), .O(n11476)
         );
  MUX2S U31719 ( .A(A67_shift[87]), .B(A67_shift[79]), .S(n13821), .O(n11475)
         );
  MUX2S U31720 ( .A(A67_shift[95]), .B(A67_shift[87]), .S(n13821), .O(n11474)
         );
  MUX2S U31721 ( .A(A67_shift[103]), .B(A67_shift[95]), .S(n13821), .O(n11473)
         );
  MUX2S U31722 ( .A(A67_shift[111]), .B(A67_shift[103]), .S(n13821), .O(n11472) );
  MUX2S U31723 ( .A(A67_shift[119]), .B(A67_shift[111]), .S(n13821), .O(n11471) );
  MUX2S U31724 ( .A(A67_shift[127]), .B(A67_shift[119]), .S(n13821), .O(n11470) );
  MUX2S U31725 ( .A(A67_shift[135]), .B(A67_shift[127]), .S(n13821), .O(n11469) );
  MUX2S U31726 ( .A(A67_shift[143]), .B(A67_shift[135]), .S(n13821), .O(n11468) );
  MUX2S U31727 ( .A(A67_shift[151]), .B(A67_shift[143]), .S(n13821), .O(n11467) );
  MUX2S U31728 ( .A(A67_shift[159]), .B(A67_shift[151]), .S(n13821), .O(n11466) );
  MUX2S U31729 ( .A(A67_shift[167]), .B(A67_shift[159]), .S(n13821), .O(n11465) );
  MUX2S U31730 ( .A(A67_shift[175]), .B(A67_shift[167]), .S(n13821), .O(n11464) );
  MUX2S U31731 ( .A(A67_shift[183]), .B(A67_shift[175]), .S(n13821), .O(n11463) );
  MUX2S U31732 ( .A(A67_shift[191]), .B(A67_shift[183]), .S(n13821), .O(n11462) );
  MUX2S U31733 ( .A(A67_shift[199]), .B(A67_shift[191]), .S(n13821), .O(n11461) );
  MUX2S U31734 ( .A(A67_shift[207]), .B(A67_shift[199]), .S(n13821), .O(n11460) );
  MUX2S U31735 ( .A(A67_shift[215]), .B(A67_shift[207]), .S(n13821), .O(n11459) );
  MUX2S U31736 ( .A(A67_shift[223]), .B(A67_shift[215]), .S(n13821), .O(n11458) );
  MUX2S U31737 ( .A(A67_shift[231]), .B(A67_shift[223]), .S(n13774), .O(n11457) );
  MUX2S U31738 ( .A(A67_shift[239]), .B(A67_shift[231]), .S(n13821), .O(n11456) );
  MUX2S U31739 ( .A(A67_shift[247]), .B(A67_shift[239]), .S(n13774), .O(n11455) );
  MUX2S U31740 ( .A(A67_shift[255]), .B(A67_shift[247]), .S(n13821), .O(n11454) );
  AOI22S U31741 ( .A1(n28412), .A2(img[15]), .B1(n24374), .B2(n31995), .O(
        n29535) );
  ND2S U31742 ( .I1(n24340), .I2(n29535), .O(n29537) );
  MUX2 U31743 ( .A(img[119]), .B(n29537), .S(n29536), .O(n13419) );
  MUX2S U31744 ( .A(rgb_value[23]), .B(image[7]), .S(in_valid), .O(n11228) );
  BUF1 U31745 ( .I(in_valid), .O(n29914) );
  MUX2S U31746 ( .A(rgb_value[15]), .B(rgb_value[23]), .S(n29914), .O(n11220)
         );
  MUX2S U31747 ( .A(rgb_value[7]), .B(rgb_value[15]), .S(n29914), .O(n11212)
         );
  MUX2S U31748 ( .A(A67_shift[209]), .B(A67_shift[201]), .S(n13774), .O(n11267) );
  MUX2S U31749 ( .A(A67_shift[217]), .B(A67_shift[209]), .S(n13821), .O(n11266) );
  MUX2S U31750 ( .A(A67_shift[225]), .B(A67_shift[217]), .S(n13774), .O(n11265) );
  MUX2S U31751 ( .A(A67_shift[233]), .B(A67_shift[225]), .S(n13821), .O(n11264) );
  MUX2S U31752 ( .A(A67_shift[241]), .B(A67_shift[233]), .S(n13774), .O(n11263) );
  MUX2S U31753 ( .A(A67_shift[249]), .B(A67_shift[241]), .S(n13821), .O(n11262) );
  NR2 U31754 ( .I1(temp_cnt[1]), .I2(temp_cnt[2]), .O(n29552) );
  INV1S U31755 ( .I(temp_cnt[3]), .O(n30025) );
  NR2 U31756 ( .I1(temp_cnt[0]), .I2(n30023), .O(n29547) );
  MUX2S U31757 ( .A(template[7]), .B(template_store[71]), .S(n29538), .O(
        n13605) );
  MUX2S U31758 ( .A(template[6]), .B(template_store[70]), .S(n29538), .O(
        n13604) );
  MUX2S U31759 ( .A(template[5]), .B(template_store[69]), .S(n29538), .O(
        n13603) );
  MUX2S U31760 ( .A(template[4]), .B(template_store[68]), .S(n29538), .O(
        n13602) );
  MUX2S U31761 ( .A(template[3]), .B(template_store[67]), .S(n29538), .O(
        n13601) );
  MUX2S U31762 ( .A(template[2]), .B(template_store[66]), .S(n29538), .O(
        n13600) );
  MUX2S U31763 ( .A(template[1]), .B(template_store[65]), .S(n29538), .O(
        n13599) );
  MUX2S U31764 ( .A(template[0]), .B(template_store[64]), .S(n29538), .O(
        n13598) );
  NR2 U31765 ( .I1(n29539), .I2(n30023), .O(n29549) );
  MUX2S U31766 ( .A(template[7]), .B(template_store[63]), .S(n29540), .O(
        n13597) );
  MUX2S U31767 ( .A(template[6]), .B(template_store[62]), .S(n29540), .O(
        n13596) );
  MUX2S U31768 ( .A(template[5]), .B(template_store[61]), .S(n29540), .O(
        n13595) );
  MUX2S U31769 ( .A(template[4]), .B(template_store[60]), .S(n29540), .O(
        n13594) );
  MUX2S U31770 ( .A(template[3]), .B(template_store[59]), .S(n29540), .O(
        n13593) );
  MUX2S U31771 ( .A(template[2]), .B(template_store[58]), .S(n29540), .O(
        n13592) );
  MUX2S U31772 ( .A(template[1]), .B(template_store[57]), .S(n29540), .O(
        n13591) );
  MUX2S U31773 ( .A(template[0]), .B(template_store[56]), .S(n29540), .O(
        n13590) );
  MUX2S U31774 ( .A(template[7]), .B(template_store[55]), .S(n29541), .O(
        n13589) );
  MUX2S U31775 ( .A(template[6]), .B(template_store[54]), .S(n29541), .O(
        n13588) );
  MUX2S U31776 ( .A(template[5]), .B(template_store[53]), .S(n29541), .O(
        n13587) );
  MUX2S U31777 ( .A(template[4]), .B(template_store[52]), .S(n29541), .O(
        n13586) );
  MUX2S U31778 ( .A(template[3]), .B(template_store[51]), .S(n29541), .O(
        n13585) );
  MUX2S U31779 ( .A(template[2]), .B(template_store[50]), .S(n29541), .O(
        n13584) );
  MUX2S U31780 ( .A(template[1]), .B(template_store[49]), .S(n29541), .O(
        n13583) );
  MUX2S U31781 ( .A(template[0]), .B(template_store[48]), .S(n29541), .O(
        n13582) );
  MUX2S U31782 ( .A(template[7]), .B(template_store[47]), .S(n29543), .O(
        n13581) );
  MUX2S U31783 ( .A(template[6]), .B(template_store[46]), .S(n29543), .O(
        n13580) );
  MUX2S U31784 ( .A(template[5]), .B(template_store[45]), .S(n29543), .O(
        n13579) );
  MUX2S U31785 ( .A(template[4]), .B(template_store[44]), .S(n29543), .O(
        n13578) );
  MUX2S U31786 ( .A(template[3]), .B(template_store[43]), .S(n29543), .O(
        n13577) );
  MUX2S U31787 ( .A(template[2]), .B(template_store[42]), .S(n29543), .O(
        n13576) );
  MUX2S U31788 ( .A(template[1]), .B(template_store[41]), .S(n29543), .O(
        n13575) );
  MUX2S U31789 ( .A(template[0]), .B(template_store[40]), .S(n29543), .O(
        n13574) );
  INV1S U31790 ( .I(temp_cnt[1]), .O(n29545) );
  MUX2S U31791 ( .A(template[7]), .B(template_store[39]), .S(n29544), .O(
        n13573) );
  MUX2S U31792 ( .A(template[6]), .B(template_store[38]), .S(n29544), .O(
        n13572) );
  MUX2S U31793 ( .A(template[5]), .B(template_store[37]), .S(n29544), .O(
        n13571) );
  MUX2S U31794 ( .A(template[4]), .B(template_store[36]), .S(n29544), .O(
        n13570) );
  MUX2S U31795 ( .A(template[3]), .B(template_store[35]), .S(n29544), .O(
        n13569) );
  MUX2S U31796 ( .A(template[2]), .B(template_store[34]), .S(n29544), .O(
        n13568) );
  MUX2S U31797 ( .A(template[1]), .B(template_store[33]), .S(n29544), .O(
        n13567) );
  MUX2S U31798 ( .A(template[0]), .B(template_store[32]), .S(n29544), .O(
        n13566) );
  MUX2S U31799 ( .A(template[7]), .B(template_store[31]), .S(n29546), .O(
        n13565) );
  MUX2S U31800 ( .A(template[6]), .B(template_store[30]), .S(n29546), .O(
        n13564) );
  MUX2S U31801 ( .A(template[5]), .B(template_store[29]), .S(n29546), .O(
        n13563) );
  MUX2S U31802 ( .A(template[4]), .B(template_store[28]), .S(n29546), .O(
        n13562) );
  MUX2S U31803 ( .A(template[3]), .B(template_store[27]), .S(n29546), .O(
        n13561) );
  MUX2S U31804 ( .A(template[2]), .B(template_store[26]), .S(n29546), .O(
        n13560) );
  MUX2S U31805 ( .A(template[1]), .B(template_store[25]), .S(n29546), .O(
        n13559) );
  MUX2S U31806 ( .A(template[0]), .B(template_store[24]), .S(n29546), .O(
        n13558) );
  MUX2S U31807 ( .A(template[7]), .B(template_store[23]), .S(n29548), .O(
        n13557) );
  MUX2S U31808 ( .A(template[6]), .B(template_store[22]), .S(n29548), .O(
        n13556) );
  MUX2S U31809 ( .A(template[5]), .B(template_store[21]), .S(n29548), .O(
        n13555) );
  MUX2S U31810 ( .A(template[4]), .B(template_store[20]), .S(n29548), .O(
        n13554) );
  MUX2S U31811 ( .A(template[3]), .B(template_store[19]), .S(n29548), .O(
        n13553) );
  MUX2S U31812 ( .A(template[2]), .B(template_store[18]), .S(n29548), .O(
        n13552) );
  MUX2S U31813 ( .A(template[1]), .B(template_store[17]), .S(n29548), .O(
        n13551) );
  MUX2S U31814 ( .A(template[0]), .B(template_store[16]), .S(n29548), .O(
        n13550) );
  MUX2S U31815 ( .A(template[7]), .B(template_store[15]), .S(n29550), .O(
        n13549) );
  MUX2S U31816 ( .A(template[6]), .B(template_store[14]), .S(n29550), .O(
        n13548) );
  MUX2S U31817 ( .A(template[5]), .B(template_store[13]), .S(n29550), .O(
        n13547) );
  MUX2S U31818 ( .A(template[4]), .B(template_store[12]), .S(n29550), .O(
        n13546) );
  MUX2S U31819 ( .A(template[3]), .B(template_store[11]), .S(n29550), .O(
        n13545) );
  MUX2S U31820 ( .A(template[2]), .B(template_store[10]), .S(n29550), .O(
        n13544) );
  MUX2S U31821 ( .A(template[1]), .B(template_store[9]), .S(n29550), .O(n13543) );
  MUX2S U31822 ( .A(template[0]), .B(template_store[8]), .S(n29550), .O(n13542) );
  NR2 U31823 ( .I1(temp_cnt[0]), .I2(n30025), .O(n29551) );
  MUX2S U31824 ( .A(template[7]), .B(template_store[7]), .S(n29553), .O(n13541) );
  MUX2S U31825 ( .A(template[6]), .B(template_store[6]), .S(n29553), .O(n13540) );
  MUX2S U31826 ( .A(template[5]), .B(template_store[5]), .S(n29553), .O(n13539) );
  MUX2S U31827 ( .A(template[4]), .B(template_store[4]), .S(n29553), .O(n13538) );
  MUX2S U31828 ( .A(template[3]), .B(template_store[3]), .S(n29553), .O(n13537) );
  MUX2S U31829 ( .A(template[2]), .B(template_store[2]), .S(n29553), .O(n13536) );
  MUX2S U31830 ( .A(template[1]), .B(template_store[1]), .S(n29553), .O(n13535) );
  MUX2S U31831 ( .A(template[0]), .B(template_store[0]), .S(n29553), .O(n13534) );
  FA1S U31832 ( .A(PE_mul[47]), .B(PE_mul[15]), .CI(PE_mul[79]), .CO(n29555), 
        .S(n29561) );
  FA1S U31833 ( .A(PE_mul[63]), .B(PE_mul[127]), .CI(PE_mul[95]), .CO(n29554), 
        .S(n29565) );
  FA1S U31834 ( .A(PE_mul[31]), .B(PE_mul[111]), .CI(PE_mul[143]), .CO(n29560), 
        .S(n29564) );
  FA1S U31835 ( .A(n29560), .B(n29559), .CI(n29558), .CO(n29556), .S(n29770)
         );
  FA1S U31836 ( .A(PE_mul[46]), .B(PE_mul[14]), .CI(PE_mul[78]), .CO(n29563), 
        .S(n29749) );
  FA1S U31837 ( .A(n29563), .B(n29562), .CI(n29561), .CO(n29558), .S(n29765)
         );
  FA1S U31838 ( .A(n29566), .B(n29565), .CI(n29564), .CO(n29771), .S(n29764)
         );
  FA1S U31839 ( .A(PE_mul[131]), .B(PE_mul[19]), .CI(PE_mul[67]), .CO(n29577), 
        .S(n29613) );
  FA1S U31840 ( .A(PE_mul[115]), .B(PE_mul[51]), .CI(PE_mul[99]), .CO(n29576), 
        .S(n29618) );
  FA1S U31841 ( .A(PE_mul[83]), .B(n29568), .CI(n29567), .CO(n29573), .S(
        n29617) );
  FA1S U31842 ( .A(PE_mul[34]), .B(PE_mul[2]), .CI(PE_mul[66]), .CO(n29567), 
        .S(n29590) );
  FA1S U31843 ( .A(n29571), .B(n29570), .CI(n29569), .CO(n29580), .S(n29627)
         );
  FA1S U31844 ( .A(n29574), .B(n29573), .CI(n29572), .CO(n29579), .S(n29626)
         );
  FA1S U31845 ( .A(PE_mul[52]), .B(PE_mul[132]), .CI(PE_mul[116]), .CO(n29589), 
        .S(n29574) );
  FA1S U31846 ( .A(PE_mul[20]), .B(PE_mul[68]), .CI(PE_mul[100]), .CO(n29588), 
        .S(n29570) );
  FA1S U31847 ( .A(PE_mul[36]), .B(PE_mul[4]), .CI(n29575), .CO(n29583), .S(
        n29571) );
  FA1S U31848 ( .A(PE_mul[84]), .B(n29577), .CI(n29576), .CO(n29581), .S(
        n29569) );
  NR2 U31849 ( .I1(n29630), .I2(n29631), .O(n29890) );
  FA1S U31850 ( .A(n29580), .B(n29579), .CI(n29578), .CO(n29632), .S(n29631)
         );
  FA1S U31851 ( .A(n29583), .B(n29582), .CI(n29581), .CO(n29638), .S(n29584)
         );
  FA1S U31852 ( .A(n29586), .B(n29585), .CI(n29584), .CO(n29637), .S(n29578)
         );
  FA1S U31853 ( .A(n29589), .B(n29588), .CI(n29587), .CO(n29644), .S(n29585)
         );
  FA1S U31854 ( .A(PE_mul[37]), .B(PE_mul[5]), .CI(PE_mul[69]), .CO(n29647), 
        .S(n29587) );
  FA1S U31855 ( .A(PE_mul[53]), .B(PE_mul[117]), .CI(PE_mul[85]), .CO(n29646), 
        .S(n29586) );
  FA1S U31856 ( .A(PE_mul[21]), .B(PE_mul[101]), .CI(PE_mul[133]), .CO(n29641), 
        .S(n29582) );
  NR2 U31857 ( .I1(n29632), .I2(n29633), .O(n29886) );
  NR2 U31858 ( .I1(n29890), .I2(n29886), .O(n29635) );
  FA1S U31859 ( .A(PE_mul[50]), .B(PE_mul[114]), .CI(PE_mul[82]), .CO(n29614), 
        .S(n29611) );
  FA1S U31860 ( .A(PE_mul[18]), .B(PE_mul[98]), .CI(PE_mul[130]), .CO(n29615), 
        .S(n29610) );
  FA1S U31861 ( .A(PE_mul[33]), .B(PE_mul[1]), .CI(PE_mul[65]), .CO(n29592), 
        .S(n29598) );
  FA1S U31862 ( .A(PE_mul[17]), .B(PE_mul[81]), .CI(PE_mul[49]), .CO(n29591), 
        .S(n29597) );
  FA1S U31863 ( .A(PE_mul[129]), .B(PE_mul[97]), .CI(PE_mul[113]), .CO(n29612), 
        .S(n29596) );
  FA1S U31864 ( .A(n29592), .B(n29591), .CI(n29590), .CO(n29616), .S(n29607)
         );
  NR2 U31865 ( .I1(n29605), .I2(n29606), .O(n29881) );
  FA1S U31866 ( .A(n29595), .B(n29594), .CI(n29593), .CO(n29609), .S(n29602)
         );
  FA1S U31867 ( .A(n29598), .B(n29597), .CI(n29596), .CO(n29608), .S(n29603)
         );
  OR2S U31868 ( .I1(n29602), .I2(n29603), .O(n29818) );
  FA1S U31869 ( .A(PE_mul[32]), .B(PE_mul[64]), .CI(PE_mul[96]), .CO(n29595), 
        .S(n29599) );
  FA1S U31870 ( .A(PE_mul[128]), .B(PE_mul[0]), .CI(PE_mul[112]), .CO(n29593), 
        .S(n29600) );
  OR2S U31871 ( .I1(n29599), .I2(n29600), .O(n29850) );
  FA1S U31872 ( .A(PE_mul[16]), .B(PE_mul[80]), .CI(PE_mul[48]), .CO(n29594), 
        .S(n29852) );
  ND2S U31873 ( .I1(n29600), .I2(n29599), .O(n29849) );
  INV1S U31874 ( .I(n29849), .O(n29601) );
  AO12S U31875 ( .B1(n29850), .B2(n29852), .A1(n29601), .O(n29820) );
  ND2S U31876 ( .I1(n29603), .I2(n29602), .O(n29817) );
  INV1S U31877 ( .I(n29817), .O(n29604) );
  AOI12HS U31878 ( .B1(n29818), .B2(n29820), .A1(n29604), .O(n29885) );
  ND2S U31879 ( .I1(n29606), .I2(n29605), .O(n29882) );
  OAI12HS U31880 ( .B1(n29881), .B2(n29885), .A1(n29882), .O(n29787) );
  FA1S U31881 ( .A(n29609), .B(n29608), .CI(n29607), .CO(n29619), .S(n29606)
         );
  FA1S U31882 ( .A(n29612), .B(n29611), .CI(n29610), .CO(n29624), .S(n29605)
         );
  FA1S U31883 ( .A(n29615), .B(n29614), .CI(n29613), .CO(n29572), .S(n29623)
         );
  FA1S U31884 ( .A(n29618), .B(n29617), .CI(n29616), .CO(n29625), .S(n29622)
         );
  OR2S U31885 ( .I1(n29619), .I2(n29620), .O(n29785) );
  ND2S U31886 ( .I1(n29620), .I2(n29619), .O(n29784) );
  INV1S U31887 ( .I(n29784), .O(n29621) );
  AOI12HS U31888 ( .B1(n29787), .B2(n29785), .A1(n29621), .O(n29857) );
  FA1S U31889 ( .A(n29624), .B(n29623), .CI(n29622), .CO(n29628), .S(n29620)
         );
  FA1S U31890 ( .A(n29627), .B(n29626), .CI(n29625), .CO(n29630), .S(n29629)
         );
  NR2 U31891 ( .I1(n29628), .I2(n29629), .O(n29853) );
  ND2S U31892 ( .I1(n29629), .I2(n29628), .O(n29854) );
  OAI12HS U31893 ( .B1(n29857), .B2(n29853), .A1(n29854), .O(n29822) );
  ND2S U31894 ( .I1(n29631), .I2(n29630), .O(n29889) );
  ND2S U31895 ( .I1(n29633), .I2(n29632), .O(n29887) );
  OAI12HS U31896 ( .B1(n29886), .B2(n29889), .A1(n29887), .O(n29634) );
  AOI12HS U31897 ( .B1(n29635), .B2(n29822), .A1(n29634), .O(n29791) );
  FA1S U31898 ( .A(n29638), .B(n29637), .CI(n29636), .CO(n29648), .S(n29633)
         );
  FA1S U31899 ( .A(n29641), .B(n29640), .CI(n29639), .CO(n29652), .S(n29642)
         );
  FA1S U31900 ( .A(n29644), .B(n29643), .CI(n29642), .CO(n29651), .S(n29636)
         );
  FA1S U31901 ( .A(n29647), .B(n29646), .CI(n29645), .CO(n29658), .S(n29643)
         );
  FA1S U31902 ( .A(PE_mul[38]), .B(PE_mul[6]), .CI(PE_mul[70]), .CO(n29661), 
        .S(n29645) );
  FA1S U31903 ( .A(PE_mul[54]), .B(PE_mul[118]), .CI(PE_mul[86]), .CO(n29660), 
        .S(n29640) );
  FA1S U31904 ( .A(PE_mul[22]), .B(PE_mul[102]), .CI(PE_mul[134]), .CO(n29655), 
        .S(n29639) );
  NR2 U31905 ( .I1(n29648), .I2(n29649), .O(n29788) );
  ND2S U31906 ( .I1(n29649), .I2(n29648), .O(n29789) );
  OAI12HS U31907 ( .B1(n29791), .B2(n29788), .A1(n29789), .O(n29862) );
  FA1S U31908 ( .A(n29652), .B(n29651), .CI(n29650), .CO(n29662), .S(n29649)
         );
  FA1S U31909 ( .A(n29655), .B(n29654), .CI(n29653), .CO(n29667), .S(n29656)
         );
  FA1S U31910 ( .A(n29658), .B(n29657), .CI(n29656), .CO(n29666), .S(n29650)
         );
  FA1S U31911 ( .A(n29661), .B(n29660), .CI(n29659), .CO(n29673), .S(n29657)
         );
  FA1S U31912 ( .A(PE_mul[39]), .B(PE_mul[7]), .CI(PE_mul[71]), .CO(n29676), 
        .S(n29659) );
  FA1S U31913 ( .A(PE_mul[55]), .B(PE_mul[119]), .CI(PE_mul[87]), .CO(n29675), 
        .S(n29654) );
  FA1S U31914 ( .A(PE_mul[23]), .B(PE_mul[103]), .CI(PE_mul[135]), .CO(n29670), 
        .S(n29653) );
  OR2S U31915 ( .I1(n29662), .I2(n29663), .O(n29861) );
  ND2S U31916 ( .I1(n29663), .I2(n29662), .O(n29860) );
  INV1S U31917 ( .I(n29860), .O(n29664) );
  AOI12HS U31918 ( .B1(n29862), .B2(n29861), .A1(n29664), .O(n29829) );
  FA1S U31919 ( .A(n29667), .B(n29666), .CI(n29665), .CO(n29677), .S(n29663)
         );
  FA1S U31920 ( .A(n29670), .B(n29669), .CI(n29668), .CO(n29681), .S(n29671)
         );
  FA1S U31921 ( .A(n29673), .B(n29672), .CI(n29671), .CO(n29680), .S(n29665)
         );
  FA1S U31922 ( .A(n29676), .B(n29675), .CI(n29674), .CO(n29687), .S(n29672)
         );
  FA1S U31923 ( .A(PE_mul[40]), .B(PE_mul[8]), .CI(PE_mul[72]), .CO(n29690), 
        .S(n29674) );
  FA1S U31924 ( .A(PE_mul[56]), .B(PE_mul[120]), .CI(PE_mul[88]), .CO(n29689), 
        .S(n29669) );
  FA1S U31925 ( .A(PE_mul[24]), .B(PE_mul[104]), .CI(PE_mul[136]), .CO(n29684), 
        .S(n29668) );
  NR2 U31926 ( .I1(n29677), .I2(n29678), .O(n29826) );
  ND2S U31927 ( .I1(n29678), .I2(n29677), .O(n29827) );
  OAI12HS U31928 ( .B1(n29829), .B2(n29826), .A1(n29827), .O(n29900) );
  FA1S U31929 ( .A(n29681), .B(n29680), .CI(n29679), .CO(n29691), .S(n29678)
         );
  FA1S U31930 ( .A(n29684), .B(n29683), .CI(n29682), .CO(n29696), .S(n29685)
         );
  FA1S U31931 ( .A(n29687), .B(n29686), .CI(n29685), .CO(n29695), .S(n29679)
         );
  FA1S U31932 ( .A(n29690), .B(n29689), .CI(n29688), .CO(n29702), .S(n29686)
         );
  FA1S U31933 ( .A(PE_mul[41]), .B(PE_mul[9]), .CI(PE_mul[73]), .CO(n29705), 
        .S(n29688) );
  FA1S U31934 ( .A(PE_mul[57]), .B(PE_mul[121]), .CI(PE_mul[89]), .CO(n29704), 
        .S(n29683) );
  FA1S U31935 ( .A(PE_mul[25]), .B(PE_mul[105]), .CI(PE_mul[137]), .CO(n29699), 
        .S(n29682) );
  OR2S U31936 ( .I1(n29691), .I2(n29692), .O(n29899) );
  ND2S U31937 ( .I1(n29692), .I2(n29691), .O(n29898) );
  INV1S U31938 ( .I(n29898), .O(n29693) );
  AOI12HS U31939 ( .B1(n29900), .B2(n29899), .A1(n29693), .O(n29799) );
  FA1S U31940 ( .A(n29696), .B(n29695), .CI(n29694), .CO(n29706), .S(n29692)
         );
  FA1S U31941 ( .A(n29699), .B(n29698), .CI(n29697), .CO(n29710), .S(n29700)
         );
  FA1S U31942 ( .A(n29702), .B(n29701), .CI(n29700), .CO(n29709), .S(n29694)
         );
  FA1S U31943 ( .A(n29705), .B(n29704), .CI(n29703), .CO(n29716), .S(n29701)
         );
  FA1S U31944 ( .A(PE_mul[42]), .B(PE_mul[10]), .CI(PE_mul[74]), .CO(n29719), 
        .S(n29703) );
  FA1S U31945 ( .A(PE_mul[58]), .B(PE_mul[122]), .CI(PE_mul[90]), .CO(n29718), 
        .S(n29698) );
  FA1S U31946 ( .A(PE_mul[26]), .B(PE_mul[106]), .CI(PE_mul[138]), .CO(n29713), 
        .S(n29697) );
  NR2 U31947 ( .I1(n29706), .I2(n29707), .O(n29796) );
  ND2S U31948 ( .I1(n29707), .I2(n29706), .O(n29797) );
  OAI12HS U31949 ( .B1(n29799), .B2(n29796), .A1(n29797), .O(n29846) );
  FA1S U31950 ( .A(n29710), .B(n29709), .CI(n29708), .CO(n29720), .S(n29707)
         );
  FA1S U31951 ( .A(n29713), .B(n29712), .CI(n29711), .CO(n29725), .S(n29714)
         );
  FA1S U31952 ( .A(n29716), .B(n29715), .CI(n29714), .CO(n29724), .S(n29708)
         );
  FA1S U31953 ( .A(n29719), .B(n29718), .CI(n29717), .CO(n29731), .S(n29715)
         );
  FA1S U31954 ( .A(PE_mul[43]), .B(PE_mul[11]), .CI(PE_mul[75]), .CO(n29734), 
        .S(n29717) );
  FA1S U31955 ( .A(PE_mul[59]), .B(PE_mul[123]), .CI(PE_mul[91]), .CO(n29733), 
        .S(n29712) );
  FA1S U31956 ( .A(PE_mul[27]), .B(PE_mul[107]), .CI(PE_mul[139]), .CO(n29728), 
        .S(n29711) );
  OR2S U31957 ( .I1(n29720), .I2(n29721), .O(n29845) );
  ND2S U31958 ( .I1(n29721), .I2(n29720), .O(n29844) );
  INV1S U31959 ( .I(n29844), .O(n29722) );
  AOI12HS U31960 ( .B1(n29846), .B2(n29845), .A1(n29722), .O(n29814) );
  FA1S U31961 ( .A(n29725), .B(n29724), .CI(n29723), .CO(n29735), .S(n29721)
         );
  FA1S U31962 ( .A(n29728), .B(n29727), .CI(n29726), .CO(n29739), .S(n29729)
         );
  FA1S U31963 ( .A(n29731), .B(n29730), .CI(n29729), .CO(n29738), .S(n29723)
         );
  FA1S U31964 ( .A(n29734), .B(n29733), .CI(n29732), .CO(n29745), .S(n29730)
         );
  FA1S U31965 ( .A(PE_mul[44]), .B(PE_mul[12]), .CI(PE_mul[76]), .CO(n29748), 
        .S(n29732) );
  FA1S U31966 ( .A(PE_mul[60]), .B(PE_mul[124]), .CI(PE_mul[92]), .CO(n29747), 
        .S(n29727) );
  FA1S U31967 ( .A(PE_mul[45]), .B(PE_mul[13]), .CI(PE_mul[77]), .CO(n29751), 
        .S(n29746) );
  FA1S U31968 ( .A(PE_mul[28]), .B(PE_mul[108]), .CI(PE_mul[140]), .CO(n29742), 
        .S(n29726) );
  FA1S U31969 ( .A(PE_mul[61]), .B(PE_mul[125]), .CI(PE_mul[93]), .CO(n29750), 
        .S(n29741) );
  NR2 U31970 ( .I1(n29735), .I2(n29736), .O(n29811) );
  ND2S U31971 ( .I1(n29736), .I2(n29735), .O(n29812) );
  OAI12HS U31972 ( .B1(n29814), .B2(n29811), .A1(n29812), .O(n29877) );
  FA1S U31973 ( .A(n29739), .B(n29738), .CI(n29737), .CO(n29752), .S(n29736)
         );
  FA1S U31974 ( .A(n29742), .B(n29741), .CI(n29740), .CO(n29757), .S(n29743)
         );
  FA1S U31975 ( .A(n29745), .B(n29744), .CI(n29743), .CO(n29756), .S(n29737)
         );
  FA1S U31976 ( .A(n29748), .B(n29747), .CI(n29746), .CO(n29763), .S(n29744)
         );
  FA1S U31977 ( .A(n29751), .B(n29750), .CI(n29749), .CO(n29766), .S(n29762)
         );
  FA1S U31978 ( .A(PE_mul[29]), .B(PE_mul[109]), .CI(PE_mul[141]), .CO(n29760), 
        .S(n29740) );
  FA1S U31979 ( .A(PE_mul[62]), .B(PE_mul[126]), .CI(PE_mul[94]), .CO(n29562), 
        .S(n29759) );
  FA1S U31980 ( .A(PE_mul[30]), .B(PE_mul[110]), .CI(PE_mul[142]), .CO(n29566), 
        .S(n29758) );
  OR2S U31981 ( .I1(n29752), .I2(n29753), .O(n29876) );
  ND2S U31982 ( .I1(n29753), .I2(n29752), .O(n29875) );
  INV1S U31983 ( .I(n29875), .O(n29754) );
  AOI12HS U31984 ( .B1(n29877), .B2(n29876), .A1(n29754), .O(n29781) );
  FA1S U31985 ( .A(n29757), .B(n29756), .CI(n29755), .CO(n29767), .S(n29753)
         );
  FA1S U31986 ( .A(n29760), .B(n29759), .CI(n29758), .CO(n29774), .S(n29761)
         );
  FA1S U31987 ( .A(n29763), .B(n29762), .CI(n29761), .CO(n29773), .S(n29755)
         );
  FA1S U31988 ( .A(n29766), .B(n29765), .CI(n29764), .CO(n29769), .S(n29772)
         );
  NR2 U31989 ( .I1(n29767), .I2(n29768), .O(n29778) );
  ND2S U31990 ( .I1(n29768), .I2(n29767), .O(n29779) );
  OAI12HS U31991 ( .B1(n29781), .B2(n29778), .A1(n29779), .O(n29842) );
  FA1S U31992 ( .A(n29771), .B(n29770), .CI(n29769), .CO(n29809), .S(n29775)
         );
  FA1S U31993 ( .A(n29774), .B(n29773), .CI(n29772), .CO(n29776), .S(n29768)
         );
  OR2S U31994 ( .I1(n29775), .I2(n29776), .O(n29841) );
  ND2S U31995 ( .I1(n29776), .I2(n29775), .O(n29840) );
  INV1S U31996 ( .I(n29840), .O(n29777) );
  INV1S U31997 ( .I(n29778), .O(n29780) );
  ND2S U31998 ( .I1(n29780), .I2(n29779), .O(n29782) );
  XOR2HS U31999 ( .I1(n29782), .I2(n29781), .O(n29783) );
  INV1S U32000 ( .I(out_cnt[3]), .O(n29801) );
  NR2 U32001 ( .I1(n29801), .I2(n29793), .O(n29879) );
  ND2S U32002 ( .I1(n29783), .I2(n29879), .O(n29805) );
  ND2S U32003 ( .I1(n29785), .I2(n29784), .O(n29786) );
  XNR2HS U32004 ( .I1(n29787), .I2(n29786), .O(n29795) );
  INV1S U32005 ( .I(n29788), .O(n29790) );
  ND2S U32006 ( .I1(n29790), .I2(n29789), .O(n29792) );
  XOR2HS U32007 ( .I1(n29792), .I2(n29791), .O(n29794) );
  NR2 U32008 ( .I1(out_cnt[3]), .I2(n29793), .O(n29894) );
  AOI22S U32009 ( .A1(n29897), .A2(n29795), .B1(n29794), .B2(n29894), .O(
        n29804) );
  INV1S U32010 ( .I(n29796), .O(n29798) );
  ND2S U32011 ( .I1(n29798), .I2(n29797), .O(n29800) );
  XOR2HS U32012 ( .I1(n29800), .I2(n29799), .O(n29802) );
  NR2 U32013 ( .I1(n29801), .I2(out_cnt[2]), .O(n29902) );
  ND2S U32014 ( .I1(n29802), .I2(n29902), .O(n29803) );
  ND3S U32015 ( .I1(n29805), .I2(n29804), .I3(n29803), .O(n29806) );
  AO12S U32016 ( .B1(n29807), .B2(out_cnt[4]), .A1(n29806), .O(n29838) );
  FA1S U32017 ( .A(n29810), .B(n29809), .CI(n29808), .CO(n29873), .S(n29836)
         );
  INV1S U32018 ( .I(n29811), .O(n29813) );
  ND2S U32019 ( .I1(n29813), .I2(n29812), .O(n29815) );
  XOR2HS U32020 ( .I1(n29815), .I2(n29814), .O(n29816) );
  ND2S U32021 ( .I1(n29816), .I2(n29879), .O(n29834) );
  ND2S U32022 ( .I1(n29818), .I2(n29817), .O(n29819) );
  XNR2HS U32023 ( .I1(n29820), .I2(n29819), .O(n29825) );
  INV1S U32024 ( .I(n29890), .O(n29821) );
  ND2S U32025 ( .I1(n29821), .I2(n29889), .O(n29823) );
  INV1S U32026 ( .I(n29822), .O(n29891) );
  XOR2HS U32027 ( .I1(n29823), .I2(n29891), .O(n29824) );
  AOI22S U32028 ( .A1(n29897), .A2(n29825), .B1(n29824), .B2(n29894), .O(
        n29833) );
  INV1S U32029 ( .I(n29826), .O(n29828) );
  ND2S U32030 ( .I1(n29828), .I2(n29827), .O(n29830) );
  XOR2HS U32031 ( .I1(n29830), .I2(n29829), .O(n29831) );
  ND2S U32032 ( .I1(n29831), .I2(n29902), .O(n29832) );
  ND3S U32033 ( .I1(n29834), .I2(n29833), .I3(n29832), .O(n29835) );
  AO12S U32034 ( .B1(n29836), .B2(out_cnt[4]), .A1(n29835), .O(n29837) );
  MUX2S U32035 ( .A(n29838), .B(n29837), .S(n30032), .O(n29839) );
  ND2S U32036 ( .I1(n29839), .I2(out_cnt[0]), .O(n29913) );
  ND2S U32037 ( .I1(n29841), .I2(n29840), .O(n29843) );
  XNR2HS U32038 ( .I1(n29843), .I2(n29842), .O(n29869) );
  ND2S U32039 ( .I1(n29845), .I2(n29844), .O(n29847) );
  XNR2HS U32040 ( .I1(n29847), .I2(n29846), .O(n29848) );
  ND2S U32041 ( .I1(n29848), .I2(n29879), .O(n29867) );
  ND2S U32042 ( .I1(n29850), .I2(n29849), .O(n29851) );
  XNR2HS U32043 ( .I1(n29852), .I2(n29851), .O(n29859) );
  INV1S U32044 ( .I(n29853), .O(n29855) );
  ND2S U32045 ( .I1(n29855), .I2(n29854), .O(n29856) );
  XOR2HS U32046 ( .I1(n29857), .I2(n29856), .O(n29858) );
  AOI22S U32047 ( .A1(n29897), .A2(n29859), .B1(n29858), .B2(n29894), .O(
        n29866) );
  ND2S U32048 ( .I1(n29861), .I2(n29860), .O(n29863) );
  XNR2HS U32049 ( .I1(n29863), .I2(n29862), .O(n29864) );
  ND2S U32050 ( .I1(n29864), .I2(n29902), .O(n29865) );
  AO12S U32051 ( .B1(n29869), .B2(out_cnt[4]), .A1(n29868), .O(n29872) );
  INV1S U32052 ( .I(n29870), .O(n29871) );
  ND2S U32053 ( .I1(n29872), .I2(n29871), .O(n29912) );
  ND2S U32054 ( .I1(n29876), .I2(n29875), .O(n29878) );
  XNR2HS U32055 ( .I1(n29878), .I2(n29877), .O(n29880) );
  ND2S U32056 ( .I1(n29880), .I2(n29879), .O(n29906) );
  INV1S U32057 ( .I(n29881), .O(n29883) );
  ND2S U32058 ( .I1(n29883), .I2(n29882), .O(n29884) );
  XOR2HS U32059 ( .I1(n29885), .I2(n29884), .O(n29896) );
  INV1S U32060 ( .I(n29886), .O(n29888) );
  ND2S U32061 ( .I1(n29888), .I2(n29887), .O(n29893) );
  OAI12HS U32062 ( .B1(n29891), .B2(n29890), .A1(n29889), .O(n29892) );
  XNR2HS U32063 ( .I1(n29893), .I2(n29892), .O(n29895) );
  AOI22S U32064 ( .A1(n29897), .A2(n29896), .B1(n29895), .B2(n29894), .O(
        n29905) );
  ND2S U32065 ( .I1(n29899), .I2(n29898), .O(n29901) );
  XNR2HS U32066 ( .I1(n29901), .I2(n29900), .O(n29903) );
  ND2S U32067 ( .I1(n29903), .I2(n29902), .O(n29904) );
  ND3S U32068 ( .I1(n29906), .I2(n29905), .I3(n29904), .O(n29907) );
  AO12S U32069 ( .B1(n29908), .B2(out_cnt[4]), .A1(n29907), .O(n29909) );
  ND3S U32070 ( .I1(n29909), .I2(out_cnt[1]), .I3(n30030), .O(n29911) );
  AOI13HS U32071 ( .B1(n29913), .B2(n29912), .B3(n29911), .A1(n29910), .O(
        N1330) );
  MUX2S U32072 ( .A(rgb_value[22]), .B(image[6]), .S(n29914), .O(n11227) );
  MUX2S U32073 ( .A(rgb_value[21]), .B(image[5]), .S(n29914), .O(n11226) );
  MUX2S U32074 ( .A(rgb_value[20]), .B(image[4]), .S(n29914), .O(n11225) );
  MUX2S U32075 ( .A(rgb_value[19]), .B(image[3]), .S(n29914), .O(n11224) );
  MUX2S U32076 ( .A(rgb_value[18]), .B(image[2]), .S(n29914), .O(n11223) );
  MUX2S U32077 ( .A(rgb_value[17]), .B(image[1]), .S(n29914), .O(n11222) );
  MUX2S U32078 ( .A(rgb_value[16]), .B(image[0]), .S(n29914), .O(n11221) );
  MUX2S U32079 ( .A(rgb_value[14]), .B(rgb_value[22]), .S(n29914), .O(n11219)
         );
  MUX2S U32080 ( .A(rgb_value[13]), .B(rgb_value[21]), .S(n29914), .O(n11218)
         );
  MUX2S U32081 ( .A(rgb_value[12]), .B(rgb_value[20]), .S(n29914), .O(n11217)
         );
  MUX2S U32082 ( .A(rgb_value[11]), .B(rgb_value[19]), .S(n29914), .O(n11216)
         );
  MUX2S U32083 ( .A(rgb_value[10]), .B(rgb_value[18]), .S(n29914), .O(n11215)
         );
  MUX2S U32084 ( .A(rgb_value[9]), .B(rgb_value[17]), .S(n29914), .O(n11214)
         );
  MUX2S U32085 ( .A(rgb_value[8]), .B(rgb_value[16]), .S(n29914), .O(n11213)
         );
  MUX2S U32086 ( .A(rgb_value[6]), .B(rgb_value[14]), .S(in_valid), .O(n11211)
         );
  MUX2S U32087 ( .A(rgb_value[5]), .B(rgb_value[13]), .S(n29914), .O(n11210)
         );
  MUX2S U32088 ( .A(rgb_value[4]), .B(rgb_value[12]), .S(n29914), .O(n11209)
         );
  MUX2S U32089 ( .A(rgb_value[3]), .B(rgb_value[11]), .S(n29914), .O(n11208)
         );
  MUX2S U32090 ( .A(rgb_value[2]), .B(rgb_value[10]), .S(n29914), .O(n11207)
         );
  MUX2S U32091 ( .A(rgb_value[1]), .B(rgb_value[9]), .S(n29914), .O(n11206) );
  MUX2S U32092 ( .A(rgb_value[0]), .B(rgb_value[8]), .S(n29914), .O(n11205) );
  XOR3S U32093 ( .I1(rgb_value[13]), .I2(rgb_value[22]), .I3(rgb_value[6]), 
        .O(intadd_8_A_4_) );
  INV1S U32094 ( .I(rgb_value[19]), .O(n29931) );
  INV1S U32095 ( .I(rgb_value[10]), .O(n29932) );
  NR2 U32096 ( .I1(n29931), .I2(n29932), .O(intadd_8_A_2_) );
  NR2 U32097 ( .I1(rgb_value[14]), .I2(rgb_value[23]), .O(n29916) );
  MOAI1S U32098 ( .A1(n29916), .A2(n29915), .B1(rgb_value[14]), .B2(
        rgb_value[23]), .O(intadd_8_B_6_) );
  XOR3S U32099 ( .I1(rgb_value[12]), .I2(rgb_value[21]), .I3(rgb_value[5]), 
        .O(intadd_8_B_3_) );
  XOR3S U32100 ( .I1(rgb_value[11]), .I2(rgb_value[20]), .I3(rgb_value[4]), 
        .O(intadd_8_B_2_) );
  XOR2HS U32101 ( .I1(rgb_value[10]), .I2(rgb_value[19]), .O(intadd_8_B_1_) );
  INV1S U32102 ( .I(rgb_value[23]), .O(n29923) );
  INV1S U32103 ( .I(rgb_value[18]), .O(n29933) );
  INV1S U32104 ( .I(rgb_value[17]), .O(n29936) );
  MUX2S U32105 ( .A(rgb_value[16]), .B(rgb_value[8]), .S(n29934), .O(n29944)
         );
  INV1S U32106 ( .I(rgb_value[14]), .O(n29924) );
  INV1S U32107 ( .I(rgb_value[9]), .O(n29935) );
  INV1S U32108 ( .I(n29945), .O(n29946) );
  INV1S U32109 ( .I(n29947), .O(n29948) );
  INV1S U32110 ( .I(n29949), .O(n29950) );
  INV1S U32111 ( .I(n29951), .O(n29952) );
  INV1S U32112 ( .I(n29953), .O(n29954) );
  INV1S U32113 ( .I(n29955), .O(n29957) );
  ND2S U32114 ( .I1(n29914), .I2(n29958), .O(n29959) );
  NR2 U32115 ( .I1(in_cnt[0]), .I2(n29959), .O(N25777) );
  NR2 U32116 ( .I1(n29960), .I2(n29959), .O(N25778) );
  MOAI1S U32117 ( .A1(act_cnt[0]), .A2(n29962), .B1(act_cnt[0]), .B2(n29961), 
        .O(n13688) );
  OAI22S U32118 ( .A1(n29966), .A2(n29965), .B1(n29964), .B2(n29963), .O(
        n13687) );
  ND2S U32119 ( .I1(n29968), .I2(n29967), .O(n29985) );
  ND2S U32120 ( .I1(cal_cnt[0]), .I2(cal_cnt[1]), .O(n29972) );
  ND2S U32121 ( .I1(n29985), .I2(n29972), .O(n29970) );
  NR2 U32122 ( .I1(n29969), .I2(n29985), .O(n29980) );
  MOAI1S U32123 ( .A1(n29971), .A2(n29970), .B1(cal_cnt[1]), .B2(n29980), .O(
        n13654) );
  INV1S U32124 ( .I(n29985), .O(n29982) );
  MOAI1S U32125 ( .A1(cal_cnt[0]), .A2(n29982), .B1(cal_cnt[0]), .B2(n29980), 
        .O(n13653) );
  MOAI1S U32126 ( .A1(n29973), .A2(n29972), .B1(n29973), .B2(n29972), .O(
        n29974) );
  MOAI1S U32127 ( .A1(n29982), .A2(n29974), .B1(cal_cnt[2]), .B2(n29980), .O(
        n13652) );
  INV1S U32128 ( .I(cal_cnt[3]), .O(n29977) );
  ND3S U32129 ( .I1(cal_cnt[0]), .I2(cal_cnt[1]), .I3(cal_cnt[2]), .O(n29976)
         );
  MOAI1S U32130 ( .A1(n29977), .A2(n29976), .B1(n29977), .B2(n29976), .O(
        n29975) );
  MOAI1S U32131 ( .A1(n29982), .A2(n29975), .B1(cal_cnt[3]), .B2(n29980), .O(
        n13651) );
  NR2 U32132 ( .I1(n29977), .I2(n29976), .O(n29979) );
  MOAI1S U32133 ( .A1(cal_cnt[4]), .A2(n29979), .B1(cal_cnt[4]), .B2(n29979), 
        .O(n29978) );
  MOAI1S U32134 ( .A1(n29982), .A2(n29978), .B1(cal_cnt[4]), .B2(n29980), .O(
        n13650) );
  INV1S U32135 ( .I(cal_cnt[5]), .O(n29984) );
  ND2S U32136 ( .I1(cal_cnt[4]), .I2(n29979), .O(n29983) );
  MOAI1S U32137 ( .A1(n29984), .A2(n29983), .B1(n29984), .B2(n29983), .O(
        n29981) );
  MOAI1S U32138 ( .A1(n29982), .A2(n29981), .B1(cal_cnt[5]), .B2(n29980), .O(
        n13649) );
  INV1S U32139 ( .I(cal_cnt[6]), .O(n29988) );
  NR2 U32140 ( .I1(n29984), .I2(n29983), .O(n29986) );
  ND2S U32141 ( .I1(n29986), .I2(n29985), .O(n29987) );
  NR2 U32142 ( .I1(n29988), .I2(n29987), .O(n29992) );
  ND2S U32143 ( .I1(n29988), .I2(n29987), .O(n29989) );
  ND2S U32144 ( .I1(n29991), .I2(n29989), .O(n29990) );
  NR2 U32145 ( .I1(n29992), .I2(n29990), .O(n13648) );
  ND2S U32146 ( .I1(cal_cnt[7]), .I2(n29992), .O(n29994) );
  AN2S U32147 ( .I1(n29991), .I2(n29994), .O(n29993) );
  OA12S U32148 ( .B1(cal_cnt[7]), .B2(n29992), .A1(n29993), .O(n13647) );
  MOAI1S U32149 ( .A1(cal_cnt[8]), .A2(n29994), .B1(cal_cnt[8]), .B2(n29993), 
        .O(n13646) );
  MOAI1S U32150 ( .A1(set_cnt[2]), .A2(n29999), .B1(n29998), .B2(n29997), .O(
        n30000) );
  MOAI1S U32151 ( .A1(set_cnt[3]), .A2(n30001), .B1(set_cnt[3]), .B2(n30000), 
        .O(n13634) );
  INV1S U32152 ( .I(addr[0]), .O(n30002) );
  MOAI1S U32153 ( .A1(n30002), .A2(n30011), .B1(n30002), .B2(n30014), .O(
        n13632) );
  ND2S U32154 ( .I1(n30005), .I2(n30014), .O(n30003) );
  OAI222S U32155 ( .A1(n30004), .A2(n30011), .B1(n30004), .B2(n30003), .C1(
        n30003), .C2(n30002), .O(n13631) );
  MOAI1S U32156 ( .A1(addr[2]), .A2(n30005), .B1(addr[2]), .B2(n30005), .O(
        n30006) );
  MOAI1S U32157 ( .A1(n30011), .A2(n30007), .B1(n30006), .B2(n30014), .O(
        n13630) );
  INV1S U32158 ( .I(n30011), .O(n30016) );
  OA12S U32159 ( .B1(addr[3]), .B2(n30008), .A1(n30012), .O(n30009) );
  AO22S U32160 ( .A1(n30016), .A2(addr[3]), .B1(n30009), .B2(n30014), .O(
        n13629) );
  INV1S U32161 ( .I(addr[4]), .O(n30013) );
  MOAI1S U32162 ( .A1(addr[4]), .A2(n30012), .B1(addr[4]), .B2(n30012), .O(
        n30010) );
  MOAI1S U32163 ( .A1(n30011), .A2(n30013), .B1(n30010), .B2(n30014), .O(
        n13628) );
  NR2 U32164 ( .I1(n30013), .I2(n30012), .O(n30015) );
  OAI12HS U32165 ( .B1(addr[5]), .B2(n30015), .A1(n30014), .O(n30017) );
  MOAI1S U32166 ( .A1(n30018), .A2(n30017), .B1(addr[5]), .B2(n30016), .O(
        n13627) );
  ND2S U32167 ( .I1(n30019), .I2(temp_cnt[0]), .O(n30020) );
  OAI22S U32168 ( .A1(n30021), .A2(n30020), .B1(n30019), .B2(temp_cnt[0]), .O(
        n13625) );
  AOI22S U32169 ( .A1(n30025), .A2(n30024), .B1(n30023), .B2(n30022), .O(
        n13622) );
  FACS1S U32170 ( .CI1(mult_x_431_n9), .B(mult_x_431_n39), .A(mult_x_431_n48), 
        .CI0(mult_x_431_n10), .CS(mult_x_431_n11), .CO1(mult_x_431_n7), .CO0(
        mult_x_431_n8), .S(PE_N57) );
  FACS1S U32171 ( .CI1(mult_x_433_n12), .B(mult_x_433_n42), .A(mult_x_433_n51), 
        .CI0(mult_x_433_n13), .CS(mult_x_433_n14), .CO1(mult_x_433_n10), .CO0(
        mult_x_433_n11), .S(PE_N89) );
  FACS1S U32172 ( .CI1(mult_x_433_n7), .B(mult_x_433_n33), .A(mult_x_433_n28), 
        .CI0(mult_x_433_n8), .CS(mult_x_433_n9), .CO1(mult_x_433_n5), .CO0(
        mult_x_433_n6), .S(PE_N91) );
  FA1S U32173 ( .A(intadd_8_B_6_), .B(rgb_value[15]), .CI(intadd_8_n2), .CO(
        intadd_8_n1), .S(gray_weight[6]) );
endmodule

