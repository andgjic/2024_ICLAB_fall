# 
#              Synchronous High Speed Single Port SRAM Compiler 
# 
#                    UMC 0.18um GenericII Logic Process
#    __________________________________________________________________________
# 
# 
#      (C) Copyright 2002-2009 Faraday Technology Corp. All Rights Reserved.
#    
#    This source code is an unpublished work belongs to Faraday Technology
#    Corp.  It is considered a trade secret and is not to be divulged or
#    used by parties who have not received written authorization from
#    Faraday Technology Corp.
#    
#    Faraday's home page can be found at:
#    http://www.faraday-tech.com/
#   
#       Module Name      : Memory_16_64
#       Words            : 64
#       Bits             : 16
#       Byte-Write       : 1
#       Aspect Ratio     : 1
#       Output Loading   : 0.05  (pf)
#       Data Slew        : 0.02  (ns)
#       CK Slew          : 0.02  (ns)
#       Power Ring Width : 2  (um)
# 
# -----------------------------------------------------------------------------
# 
#       Library          : FSA0M_A
#       Memaker          : 200901.2.1
#       Date             : 2024/10/27 12:34:50
# 
# -----------------------------------------------------------------------------


NAMESCASESENSITIVE ON ;
MACRO Memory_16_64
CLASS BLOCK ;
FOREIGN Memory_16_64 0.000 0.000 ;
ORIGIN 0.000 0.000 ;
SIZE 305.660 BY 156.800 ;
SYMMETRY x y r90 ;
SITE core ;
PIN GND
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
 PORT
  LAYER ME4 ;
  RECT 304.540 129.700 305.660 132.940 ;
  LAYER ME3 ;
  RECT 304.540 129.700 305.660 132.940 ;
  LAYER ME2 ;
  RECT 304.540 129.700 305.660 132.940 ;
  LAYER ME1 ;
  RECT 304.540 129.700 305.660 132.940 ;
 END
 PORT
  LAYER ME4 ;
  RECT 304.540 121.860 305.660 125.100 ;
  LAYER ME3 ;
  RECT 304.540 121.860 305.660 125.100 ;
  LAYER ME2 ;
  RECT 304.540 121.860 305.660 125.100 ;
  LAYER ME1 ;
  RECT 304.540 121.860 305.660 125.100 ;
 END
 PORT
  LAYER ME4 ;
  RECT 304.540 114.020 305.660 117.260 ;
  LAYER ME3 ;
  RECT 304.540 114.020 305.660 117.260 ;
  LAYER ME2 ;
  RECT 304.540 114.020 305.660 117.260 ;
  LAYER ME1 ;
  RECT 304.540 114.020 305.660 117.260 ;
 END
 PORT
  LAYER ME4 ;
  RECT 304.540 106.180 305.660 109.420 ;
  LAYER ME3 ;
  RECT 304.540 106.180 305.660 109.420 ;
  LAYER ME2 ;
  RECT 304.540 106.180 305.660 109.420 ;
  LAYER ME1 ;
  RECT 304.540 106.180 305.660 109.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 304.540 98.340 305.660 101.580 ;
  LAYER ME3 ;
  RECT 304.540 98.340 305.660 101.580 ;
  LAYER ME2 ;
  RECT 304.540 98.340 305.660 101.580 ;
  LAYER ME1 ;
  RECT 304.540 98.340 305.660 101.580 ;
 END
 PORT
  LAYER ME4 ;
  RECT 304.540 90.500 305.660 93.740 ;
  LAYER ME3 ;
  RECT 304.540 90.500 305.660 93.740 ;
  LAYER ME2 ;
  RECT 304.540 90.500 305.660 93.740 ;
  LAYER ME1 ;
  RECT 304.540 90.500 305.660 93.740 ;
 END
 PORT
  LAYER ME4 ;
  RECT 304.540 51.300 305.660 54.540 ;
  LAYER ME3 ;
  RECT 304.540 51.300 305.660 54.540 ;
  LAYER ME2 ;
  RECT 304.540 51.300 305.660 54.540 ;
  LAYER ME1 ;
  RECT 304.540 51.300 305.660 54.540 ;
 END
 PORT
  LAYER ME4 ;
  RECT 304.540 43.460 305.660 46.700 ;
  LAYER ME3 ;
  RECT 304.540 43.460 305.660 46.700 ;
  LAYER ME2 ;
  RECT 304.540 43.460 305.660 46.700 ;
  LAYER ME1 ;
  RECT 304.540 43.460 305.660 46.700 ;
 END
 PORT
  LAYER ME4 ;
  RECT 304.540 35.620 305.660 38.860 ;
  LAYER ME3 ;
  RECT 304.540 35.620 305.660 38.860 ;
  LAYER ME2 ;
  RECT 304.540 35.620 305.660 38.860 ;
  LAYER ME1 ;
  RECT 304.540 35.620 305.660 38.860 ;
 END
 PORT
  LAYER ME4 ;
  RECT 304.540 27.780 305.660 31.020 ;
  LAYER ME3 ;
  RECT 304.540 27.780 305.660 31.020 ;
  LAYER ME2 ;
  RECT 304.540 27.780 305.660 31.020 ;
  LAYER ME1 ;
  RECT 304.540 27.780 305.660 31.020 ;
 END
 PORT
  LAYER ME4 ;
  RECT 304.540 19.940 305.660 23.180 ;
  LAYER ME3 ;
  RECT 304.540 19.940 305.660 23.180 ;
  LAYER ME2 ;
  RECT 304.540 19.940 305.660 23.180 ;
  LAYER ME1 ;
  RECT 304.540 19.940 305.660 23.180 ;
 END
 PORT
  LAYER ME4 ;
  RECT 304.540 12.100 305.660 15.340 ;
  LAYER ME3 ;
  RECT 304.540 12.100 305.660 15.340 ;
  LAYER ME2 ;
  RECT 304.540 12.100 305.660 15.340 ;
  LAYER ME1 ;
  RECT 304.540 12.100 305.660 15.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 129.700 1.120 132.940 ;
  LAYER ME3 ;
  RECT 0.000 129.700 1.120 132.940 ;
  LAYER ME2 ;
  RECT 0.000 129.700 1.120 132.940 ;
  LAYER ME1 ;
  RECT 0.000 129.700 1.120 132.940 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 121.860 1.120 125.100 ;
  LAYER ME3 ;
  RECT 0.000 121.860 1.120 125.100 ;
  LAYER ME2 ;
  RECT 0.000 121.860 1.120 125.100 ;
  LAYER ME1 ;
  RECT 0.000 121.860 1.120 125.100 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 114.020 1.120 117.260 ;
  LAYER ME3 ;
  RECT 0.000 114.020 1.120 117.260 ;
  LAYER ME2 ;
  RECT 0.000 114.020 1.120 117.260 ;
  LAYER ME1 ;
  RECT 0.000 114.020 1.120 117.260 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 106.180 1.120 109.420 ;
  LAYER ME3 ;
  RECT 0.000 106.180 1.120 109.420 ;
  LAYER ME2 ;
  RECT 0.000 106.180 1.120 109.420 ;
  LAYER ME1 ;
  RECT 0.000 106.180 1.120 109.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 98.340 1.120 101.580 ;
  LAYER ME3 ;
  RECT 0.000 98.340 1.120 101.580 ;
  LAYER ME2 ;
  RECT 0.000 98.340 1.120 101.580 ;
  LAYER ME1 ;
  RECT 0.000 98.340 1.120 101.580 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 90.500 1.120 93.740 ;
  LAYER ME3 ;
  RECT 0.000 90.500 1.120 93.740 ;
  LAYER ME2 ;
  RECT 0.000 90.500 1.120 93.740 ;
  LAYER ME1 ;
  RECT 0.000 90.500 1.120 93.740 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 51.300 1.120 54.540 ;
  LAYER ME3 ;
  RECT 0.000 51.300 1.120 54.540 ;
  LAYER ME2 ;
  RECT 0.000 51.300 1.120 54.540 ;
  LAYER ME1 ;
  RECT 0.000 51.300 1.120 54.540 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 43.460 1.120 46.700 ;
  LAYER ME3 ;
  RECT 0.000 43.460 1.120 46.700 ;
  LAYER ME2 ;
  RECT 0.000 43.460 1.120 46.700 ;
  LAYER ME1 ;
  RECT 0.000 43.460 1.120 46.700 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 35.620 1.120 38.860 ;
  LAYER ME3 ;
  RECT 0.000 35.620 1.120 38.860 ;
  LAYER ME2 ;
  RECT 0.000 35.620 1.120 38.860 ;
  LAYER ME1 ;
  RECT 0.000 35.620 1.120 38.860 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 27.780 1.120 31.020 ;
  LAYER ME3 ;
  RECT 0.000 27.780 1.120 31.020 ;
  LAYER ME2 ;
  RECT 0.000 27.780 1.120 31.020 ;
  LAYER ME1 ;
  RECT 0.000 27.780 1.120 31.020 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 19.940 1.120 23.180 ;
  LAYER ME3 ;
  RECT 0.000 19.940 1.120 23.180 ;
  LAYER ME2 ;
  RECT 0.000 19.940 1.120 23.180 ;
  LAYER ME1 ;
  RECT 0.000 19.940 1.120 23.180 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 12.100 1.120 15.340 ;
  LAYER ME3 ;
  RECT 0.000 12.100 1.120 15.340 ;
  LAYER ME2 ;
  RECT 0.000 12.100 1.120 15.340 ;
  LAYER ME1 ;
  RECT 0.000 12.100 1.120 15.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 289.940 155.680 293.480 156.800 ;
  LAYER ME3 ;
  RECT 289.940 155.680 293.480 156.800 ;
  LAYER ME2 ;
  RECT 289.940 155.680 293.480 156.800 ;
  LAYER ME1 ;
  RECT 289.940 155.680 293.480 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 281.260 155.680 284.800 156.800 ;
  LAYER ME3 ;
  RECT 281.260 155.680 284.800 156.800 ;
  LAYER ME2 ;
  RECT 281.260 155.680 284.800 156.800 ;
  LAYER ME1 ;
  RECT 281.260 155.680 284.800 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 272.580 155.680 276.120 156.800 ;
  LAYER ME3 ;
  RECT 272.580 155.680 276.120 156.800 ;
  LAYER ME2 ;
  RECT 272.580 155.680 276.120 156.800 ;
  LAYER ME1 ;
  RECT 272.580 155.680 276.120 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 229.180 155.680 232.720 156.800 ;
  LAYER ME3 ;
  RECT 229.180 155.680 232.720 156.800 ;
  LAYER ME2 ;
  RECT 229.180 155.680 232.720 156.800 ;
  LAYER ME1 ;
  RECT 229.180 155.680 232.720 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 220.500 155.680 224.040 156.800 ;
  LAYER ME3 ;
  RECT 220.500 155.680 224.040 156.800 ;
  LAYER ME2 ;
  RECT 220.500 155.680 224.040 156.800 ;
  LAYER ME1 ;
  RECT 220.500 155.680 224.040 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 211.820 155.680 215.360 156.800 ;
  LAYER ME3 ;
  RECT 211.820 155.680 215.360 156.800 ;
  LAYER ME2 ;
  RECT 211.820 155.680 215.360 156.800 ;
  LAYER ME1 ;
  RECT 211.820 155.680 215.360 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 203.140 155.680 206.680 156.800 ;
  LAYER ME3 ;
  RECT 203.140 155.680 206.680 156.800 ;
  LAYER ME2 ;
  RECT 203.140 155.680 206.680 156.800 ;
  LAYER ME1 ;
  RECT 203.140 155.680 206.680 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 194.460 155.680 198.000 156.800 ;
  LAYER ME3 ;
  RECT 194.460 155.680 198.000 156.800 ;
  LAYER ME2 ;
  RECT 194.460 155.680 198.000 156.800 ;
  LAYER ME1 ;
  RECT 194.460 155.680 198.000 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 185.780 155.680 189.320 156.800 ;
  LAYER ME3 ;
  RECT 185.780 155.680 189.320 156.800 ;
  LAYER ME2 ;
  RECT 185.780 155.680 189.320 156.800 ;
  LAYER ME1 ;
  RECT 185.780 155.680 189.320 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 142.380 155.680 145.920 156.800 ;
  LAYER ME3 ;
  RECT 142.380 155.680 145.920 156.800 ;
  LAYER ME2 ;
  RECT 142.380 155.680 145.920 156.800 ;
  LAYER ME1 ;
  RECT 142.380 155.680 145.920 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 133.700 155.680 137.240 156.800 ;
  LAYER ME3 ;
  RECT 133.700 155.680 137.240 156.800 ;
  LAYER ME2 ;
  RECT 133.700 155.680 137.240 156.800 ;
  LAYER ME1 ;
  RECT 133.700 155.680 137.240 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 125.020 155.680 128.560 156.800 ;
  LAYER ME3 ;
  RECT 125.020 155.680 128.560 156.800 ;
  LAYER ME2 ;
  RECT 125.020 155.680 128.560 156.800 ;
  LAYER ME1 ;
  RECT 125.020 155.680 128.560 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 116.340 155.680 119.880 156.800 ;
  LAYER ME3 ;
  RECT 116.340 155.680 119.880 156.800 ;
  LAYER ME2 ;
  RECT 116.340 155.680 119.880 156.800 ;
  LAYER ME1 ;
  RECT 116.340 155.680 119.880 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 107.660 155.680 111.200 156.800 ;
  LAYER ME3 ;
  RECT 107.660 155.680 111.200 156.800 ;
  LAYER ME2 ;
  RECT 107.660 155.680 111.200 156.800 ;
  LAYER ME1 ;
  RECT 107.660 155.680 111.200 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 98.980 155.680 102.520 156.800 ;
  LAYER ME3 ;
  RECT 98.980 155.680 102.520 156.800 ;
  LAYER ME2 ;
  RECT 98.980 155.680 102.520 156.800 ;
  LAYER ME1 ;
  RECT 98.980 155.680 102.520 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 55.580 155.680 59.120 156.800 ;
  LAYER ME3 ;
  RECT 55.580 155.680 59.120 156.800 ;
  LAYER ME2 ;
  RECT 55.580 155.680 59.120 156.800 ;
  LAYER ME1 ;
  RECT 55.580 155.680 59.120 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 46.900 155.680 50.440 156.800 ;
  LAYER ME3 ;
  RECT 46.900 155.680 50.440 156.800 ;
  LAYER ME2 ;
  RECT 46.900 155.680 50.440 156.800 ;
  LAYER ME1 ;
  RECT 46.900 155.680 50.440 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 38.220 155.680 41.760 156.800 ;
  LAYER ME3 ;
  RECT 38.220 155.680 41.760 156.800 ;
  LAYER ME2 ;
  RECT 38.220 155.680 41.760 156.800 ;
  LAYER ME1 ;
  RECT 38.220 155.680 41.760 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 29.540 155.680 33.080 156.800 ;
  LAYER ME3 ;
  RECT 29.540 155.680 33.080 156.800 ;
  LAYER ME2 ;
  RECT 29.540 155.680 33.080 156.800 ;
  LAYER ME1 ;
  RECT 29.540 155.680 33.080 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 20.860 155.680 24.400 156.800 ;
  LAYER ME3 ;
  RECT 20.860 155.680 24.400 156.800 ;
  LAYER ME2 ;
  RECT 20.860 155.680 24.400 156.800 ;
  LAYER ME1 ;
  RECT 20.860 155.680 24.400 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 12.180 155.680 15.720 156.800 ;
  LAYER ME3 ;
  RECT 12.180 155.680 15.720 156.800 ;
  LAYER ME2 ;
  RECT 12.180 155.680 15.720 156.800 ;
  LAYER ME1 ;
  RECT 12.180 155.680 15.720 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 286.220 0.000 289.760 1.120 ;
  LAYER ME3 ;
  RECT 286.220 0.000 289.760 1.120 ;
  LAYER ME2 ;
  RECT 286.220 0.000 289.760 1.120 ;
  LAYER ME1 ;
  RECT 286.220 0.000 289.760 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 264.520 0.000 268.060 1.120 ;
  LAYER ME3 ;
  RECT 264.520 0.000 268.060 1.120 ;
  LAYER ME2 ;
  RECT 264.520 0.000 268.060 1.120 ;
  LAYER ME1 ;
  RECT 264.520 0.000 268.060 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 242.820 0.000 246.360 1.120 ;
  LAYER ME3 ;
  RECT 242.820 0.000 246.360 1.120 ;
  LAYER ME2 ;
  RECT 242.820 0.000 246.360 1.120 ;
  LAYER ME1 ;
  RECT 242.820 0.000 246.360 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 133.080 0.000 136.620 1.120 ;
  LAYER ME3 ;
  RECT 133.080 0.000 136.620 1.120 ;
  LAYER ME2 ;
  RECT 133.080 0.000 136.620 1.120 ;
  LAYER ME1 ;
  RECT 133.080 0.000 136.620 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 113.860 0.000 117.400 1.120 ;
  LAYER ME3 ;
  RECT 113.860 0.000 117.400 1.120 ;
  LAYER ME2 ;
  RECT 113.860 0.000 117.400 1.120 ;
  LAYER ME1 ;
  RECT 113.860 0.000 117.400 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 92.160 0.000 95.700 1.120 ;
  LAYER ME3 ;
  RECT 92.160 0.000 95.700 1.120 ;
  LAYER ME2 ;
  RECT 92.160 0.000 95.700 1.120 ;
  LAYER ME1 ;
  RECT 92.160 0.000 95.700 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 70.460 0.000 74.000 1.120 ;
  LAYER ME3 ;
  RECT 70.460 0.000 74.000 1.120 ;
  LAYER ME2 ;
  RECT 70.460 0.000 74.000 1.120 ;
  LAYER ME1 ;
  RECT 70.460 0.000 74.000 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 43.800 0.000 47.340 1.120 ;
  LAYER ME3 ;
  RECT 43.800 0.000 47.340 1.120 ;
  LAYER ME2 ;
  RECT 43.800 0.000 47.340 1.120 ;
  LAYER ME1 ;
  RECT 43.800 0.000 47.340 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 27.060 0.000 30.600 1.120 ;
  LAYER ME3 ;
  RECT 27.060 0.000 30.600 1.120 ;
  LAYER ME2 ;
  RECT 27.060 0.000 30.600 1.120 ;
  LAYER ME1 ;
  RECT 27.060 0.000 30.600 1.120 ;
 END
END GND
PIN VCC
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
 PORT
  LAYER ME4 ;
  RECT 304.540 125.780 305.660 129.020 ;
  LAYER ME3 ;
  RECT 304.540 125.780 305.660 129.020 ;
  LAYER ME2 ;
  RECT 304.540 125.780 305.660 129.020 ;
  LAYER ME1 ;
  RECT 304.540 125.780 305.660 129.020 ;
 END
 PORT
  LAYER ME4 ;
  RECT 304.540 117.940 305.660 121.180 ;
  LAYER ME3 ;
  RECT 304.540 117.940 305.660 121.180 ;
  LAYER ME2 ;
  RECT 304.540 117.940 305.660 121.180 ;
  LAYER ME1 ;
  RECT 304.540 117.940 305.660 121.180 ;
 END
 PORT
  LAYER ME4 ;
  RECT 304.540 110.100 305.660 113.340 ;
  LAYER ME3 ;
  RECT 304.540 110.100 305.660 113.340 ;
  LAYER ME2 ;
  RECT 304.540 110.100 305.660 113.340 ;
  LAYER ME1 ;
  RECT 304.540 110.100 305.660 113.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 304.540 102.260 305.660 105.500 ;
  LAYER ME3 ;
  RECT 304.540 102.260 305.660 105.500 ;
  LAYER ME2 ;
  RECT 304.540 102.260 305.660 105.500 ;
  LAYER ME1 ;
  RECT 304.540 102.260 305.660 105.500 ;
 END
 PORT
  LAYER ME4 ;
  RECT 304.540 94.420 305.660 97.660 ;
  LAYER ME3 ;
  RECT 304.540 94.420 305.660 97.660 ;
  LAYER ME2 ;
  RECT 304.540 94.420 305.660 97.660 ;
  LAYER ME1 ;
  RECT 304.540 94.420 305.660 97.660 ;
 END
 PORT
  LAYER ME4 ;
  RECT 304.540 86.580 305.660 89.820 ;
  LAYER ME3 ;
  RECT 304.540 86.580 305.660 89.820 ;
  LAYER ME2 ;
  RECT 304.540 86.580 305.660 89.820 ;
  LAYER ME1 ;
  RECT 304.540 86.580 305.660 89.820 ;
 END
 PORT
  LAYER ME4 ;
  RECT 304.540 47.380 305.660 50.620 ;
  LAYER ME3 ;
  RECT 304.540 47.380 305.660 50.620 ;
  LAYER ME2 ;
  RECT 304.540 47.380 305.660 50.620 ;
  LAYER ME1 ;
  RECT 304.540 47.380 305.660 50.620 ;
 END
 PORT
  LAYER ME4 ;
  RECT 304.540 39.540 305.660 42.780 ;
  LAYER ME3 ;
  RECT 304.540 39.540 305.660 42.780 ;
  LAYER ME2 ;
  RECT 304.540 39.540 305.660 42.780 ;
  LAYER ME1 ;
  RECT 304.540 39.540 305.660 42.780 ;
 END
 PORT
  LAYER ME4 ;
  RECT 304.540 31.700 305.660 34.940 ;
  LAYER ME3 ;
  RECT 304.540 31.700 305.660 34.940 ;
  LAYER ME2 ;
  RECT 304.540 31.700 305.660 34.940 ;
  LAYER ME1 ;
  RECT 304.540 31.700 305.660 34.940 ;
 END
 PORT
  LAYER ME4 ;
  RECT 304.540 23.860 305.660 27.100 ;
  LAYER ME3 ;
  RECT 304.540 23.860 305.660 27.100 ;
  LAYER ME2 ;
  RECT 304.540 23.860 305.660 27.100 ;
  LAYER ME1 ;
  RECT 304.540 23.860 305.660 27.100 ;
 END
 PORT
  LAYER ME4 ;
  RECT 304.540 16.020 305.660 19.260 ;
  LAYER ME3 ;
  RECT 304.540 16.020 305.660 19.260 ;
  LAYER ME2 ;
  RECT 304.540 16.020 305.660 19.260 ;
  LAYER ME1 ;
  RECT 304.540 16.020 305.660 19.260 ;
 END
 PORT
  LAYER ME4 ;
  RECT 304.540 8.180 305.660 11.420 ;
  LAYER ME3 ;
  RECT 304.540 8.180 305.660 11.420 ;
  LAYER ME2 ;
  RECT 304.540 8.180 305.660 11.420 ;
  LAYER ME1 ;
  RECT 304.540 8.180 305.660 11.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 125.780 1.120 129.020 ;
  LAYER ME3 ;
  RECT 0.000 125.780 1.120 129.020 ;
  LAYER ME2 ;
  RECT 0.000 125.780 1.120 129.020 ;
  LAYER ME1 ;
  RECT 0.000 125.780 1.120 129.020 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 117.940 1.120 121.180 ;
  LAYER ME3 ;
  RECT 0.000 117.940 1.120 121.180 ;
  LAYER ME2 ;
  RECT 0.000 117.940 1.120 121.180 ;
  LAYER ME1 ;
  RECT 0.000 117.940 1.120 121.180 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 110.100 1.120 113.340 ;
  LAYER ME3 ;
  RECT 0.000 110.100 1.120 113.340 ;
  LAYER ME2 ;
  RECT 0.000 110.100 1.120 113.340 ;
  LAYER ME1 ;
  RECT 0.000 110.100 1.120 113.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 102.260 1.120 105.500 ;
  LAYER ME3 ;
  RECT 0.000 102.260 1.120 105.500 ;
  LAYER ME2 ;
  RECT 0.000 102.260 1.120 105.500 ;
  LAYER ME1 ;
  RECT 0.000 102.260 1.120 105.500 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 94.420 1.120 97.660 ;
  LAYER ME3 ;
  RECT 0.000 94.420 1.120 97.660 ;
  LAYER ME2 ;
  RECT 0.000 94.420 1.120 97.660 ;
  LAYER ME1 ;
  RECT 0.000 94.420 1.120 97.660 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 86.580 1.120 89.820 ;
  LAYER ME3 ;
  RECT 0.000 86.580 1.120 89.820 ;
  LAYER ME2 ;
  RECT 0.000 86.580 1.120 89.820 ;
  LAYER ME1 ;
  RECT 0.000 86.580 1.120 89.820 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 47.380 1.120 50.620 ;
  LAYER ME3 ;
  RECT 0.000 47.380 1.120 50.620 ;
  LAYER ME2 ;
  RECT 0.000 47.380 1.120 50.620 ;
  LAYER ME1 ;
  RECT 0.000 47.380 1.120 50.620 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 39.540 1.120 42.780 ;
  LAYER ME3 ;
  RECT 0.000 39.540 1.120 42.780 ;
  LAYER ME2 ;
  RECT 0.000 39.540 1.120 42.780 ;
  LAYER ME1 ;
  RECT 0.000 39.540 1.120 42.780 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 31.700 1.120 34.940 ;
  LAYER ME3 ;
  RECT 0.000 31.700 1.120 34.940 ;
  LAYER ME2 ;
  RECT 0.000 31.700 1.120 34.940 ;
  LAYER ME1 ;
  RECT 0.000 31.700 1.120 34.940 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 23.860 1.120 27.100 ;
  LAYER ME3 ;
  RECT 0.000 23.860 1.120 27.100 ;
  LAYER ME2 ;
  RECT 0.000 23.860 1.120 27.100 ;
  LAYER ME1 ;
  RECT 0.000 23.860 1.120 27.100 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 16.020 1.120 19.260 ;
  LAYER ME3 ;
  RECT 0.000 16.020 1.120 19.260 ;
  LAYER ME2 ;
  RECT 0.000 16.020 1.120 19.260 ;
  LAYER ME1 ;
  RECT 0.000 16.020 1.120 19.260 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 8.180 1.120 11.420 ;
  LAYER ME3 ;
  RECT 0.000 8.180 1.120 11.420 ;
  LAYER ME2 ;
  RECT 0.000 8.180 1.120 11.420 ;
  LAYER ME1 ;
  RECT 0.000 8.180 1.120 11.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 294.280 155.680 297.820 156.800 ;
  LAYER ME3 ;
  RECT 294.280 155.680 297.820 156.800 ;
  LAYER ME2 ;
  RECT 294.280 155.680 297.820 156.800 ;
  LAYER ME1 ;
  RECT 294.280 155.680 297.820 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 285.600 155.680 289.140 156.800 ;
  LAYER ME3 ;
  RECT 285.600 155.680 289.140 156.800 ;
  LAYER ME2 ;
  RECT 285.600 155.680 289.140 156.800 ;
  LAYER ME1 ;
  RECT 285.600 155.680 289.140 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 276.920 155.680 280.460 156.800 ;
  LAYER ME3 ;
  RECT 276.920 155.680 280.460 156.800 ;
  LAYER ME2 ;
  RECT 276.920 155.680 280.460 156.800 ;
  LAYER ME1 ;
  RECT 276.920 155.680 280.460 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 268.240 155.680 271.780 156.800 ;
  LAYER ME3 ;
  RECT 268.240 155.680 271.780 156.800 ;
  LAYER ME2 ;
  RECT 268.240 155.680 271.780 156.800 ;
  LAYER ME1 ;
  RECT 268.240 155.680 271.780 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 224.840 155.680 228.380 156.800 ;
  LAYER ME3 ;
  RECT 224.840 155.680 228.380 156.800 ;
  LAYER ME2 ;
  RECT 224.840 155.680 228.380 156.800 ;
  LAYER ME1 ;
  RECT 224.840 155.680 228.380 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 216.160 155.680 219.700 156.800 ;
  LAYER ME3 ;
  RECT 216.160 155.680 219.700 156.800 ;
  LAYER ME2 ;
  RECT 216.160 155.680 219.700 156.800 ;
  LAYER ME1 ;
  RECT 216.160 155.680 219.700 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 207.480 155.680 211.020 156.800 ;
  LAYER ME3 ;
  RECT 207.480 155.680 211.020 156.800 ;
  LAYER ME2 ;
  RECT 207.480 155.680 211.020 156.800 ;
  LAYER ME1 ;
  RECT 207.480 155.680 211.020 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 198.800 155.680 202.340 156.800 ;
  LAYER ME3 ;
  RECT 198.800 155.680 202.340 156.800 ;
  LAYER ME2 ;
  RECT 198.800 155.680 202.340 156.800 ;
  LAYER ME1 ;
  RECT 198.800 155.680 202.340 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 190.120 155.680 193.660 156.800 ;
  LAYER ME3 ;
  RECT 190.120 155.680 193.660 156.800 ;
  LAYER ME2 ;
  RECT 190.120 155.680 193.660 156.800 ;
  LAYER ME1 ;
  RECT 190.120 155.680 193.660 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 181.440 155.680 184.980 156.800 ;
  LAYER ME3 ;
  RECT 181.440 155.680 184.980 156.800 ;
  LAYER ME2 ;
  RECT 181.440 155.680 184.980 156.800 ;
  LAYER ME1 ;
  RECT 181.440 155.680 184.980 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 138.040 155.680 141.580 156.800 ;
  LAYER ME3 ;
  RECT 138.040 155.680 141.580 156.800 ;
  LAYER ME2 ;
  RECT 138.040 155.680 141.580 156.800 ;
  LAYER ME1 ;
  RECT 138.040 155.680 141.580 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 129.360 155.680 132.900 156.800 ;
  LAYER ME3 ;
  RECT 129.360 155.680 132.900 156.800 ;
  LAYER ME2 ;
  RECT 129.360 155.680 132.900 156.800 ;
  LAYER ME1 ;
  RECT 129.360 155.680 132.900 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 120.680 155.680 124.220 156.800 ;
  LAYER ME3 ;
  RECT 120.680 155.680 124.220 156.800 ;
  LAYER ME2 ;
  RECT 120.680 155.680 124.220 156.800 ;
  LAYER ME1 ;
  RECT 120.680 155.680 124.220 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 112.000 155.680 115.540 156.800 ;
  LAYER ME3 ;
  RECT 112.000 155.680 115.540 156.800 ;
  LAYER ME2 ;
  RECT 112.000 155.680 115.540 156.800 ;
  LAYER ME1 ;
  RECT 112.000 155.680 115.540 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 103.320 155.680 106.860 156.800 ;
  LAYER ME3 ;
  RECT 103.320 155.680 106.860 156.800 ;
  LAYER ME2 ;
  RECT 103.320 155.680 106.860 156.800 ;
  LAYER ME1 ;
  RECT 103.320 155.680 106.860 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 94.640 155.680 98.180 156.800 ;
  LAYER ME3 ;
  RECT 94.640 155.680 98.180 156.800 ;
  LAYER ME2 ;
  RECT 94.640 155.680 98.180 156.800 ;
  LAYER ME1 ;
  RECT 94.640 155.680 98.180 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 51.240 155.680 54.780 156.800 ;
  LAYER ME3 ;
  RECT 51.240 155.680 54.780 156.800 ;
  LAYER ME2 ;
  RECT 51.240 155.680 54.780 156.800 ;
  LAYER ME1 ;
  RECT 51.240 155.680 54.780 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 42.560 155.680 46.100 156.800 ;
  LAYER ME3 ;
  RECT 42.560 155.680 46.100 156.800 ;
  LAYER ME2 ;
  RECT 42.560 155.680 46.100 156.800 ;
  LAYER ME1 ;
  RECT 42.560 155.680 46.100 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 33.880 155.680 37.420 156.800 ;
  LAYER ME3 ;
  RECT 33.880 155.680 37.420 156.800 ;
  LAYER ME2 ;
  RECT 33.880 155.680 37.420 156.800 ;
  LAYER ME1 ;
  RECT 33.880 155.680 37.420 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 25.200 155.680 28.740 156.800 ;
  LAYER ME3 ;
  RECT 25.200 155.680 28.740 156.800 ;
  LAYER ME2 ;
  RECT 25.200 155.680 28.740 156.800 ;
  LAYER ME1 ;
  RECT 25.200 155.680 28.740 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 16.520 155.680 20.060 156.800 ;
  LAYER ME3 ;
  RECT 16.520 155.680 20.060 156.800 ;
  LAYER ME2 ;
  RECT 16.520 155.680 20.060 156.800 ;
  LAYER ME1 ;
  RECT 16.520 155.680 20.060 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 7.840 155.680 11.380 156.800 ;
  LAYER ME3 ;
  RECT 7.840 155.680 11.380 156.800 ;
  LAYER ME2 ;
  RECT 7.840 155.680 11.380 156.800 ;
  LAYER ME1 ;
  RECT 7.840 155.680 11.380 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 294.280 0.000 297.820 1.120 ;
  LAYER ME3 ;
  RECT 294.280 0.000 297.820 1.120 ;
  LAYER ME2 ;
  RECT 294.280 0.000 297.820 1.120 ;
  LAYER ME1 ;
  RECT 294.280 0.000 297.820 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 272.580 0.000 276.120 1.120 ;
  LAYER ME3 ;
  RECT 272.580 0.000 276.120 1.120 ;
  LAYER ME2 ;
  RECT 272.580 0.000 276.120 1.120 ;
  LAYER ME1 ;
  RECT 272.580 0.000 276.120 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 255.840 0.000 259.380 1.120 ;
  LAYER ME3 ;
  RECT 255.840 0.000 259.380 1.120 ;
  LAYER ME2 ;
  RECT 255.840 0.000 259.380 1.120 ;
  LAYER ME1 ;
  RECT 255.840 0.000 259.380 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 229.180 0.000 232.720 1.120 ;
  LAYER ME3 ;
  RECT 229.180 0.000 232.720 1.120 ;
  LAYER ME2 ;
  RECT 229.180 0.000 232.720 1.120 ;
  LAYER ME1 ;
  RECT 229.180 0.000 232.720 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 121.920 0.000 125.460 1.120 ;
  LAYER ME3 ;
  RECT 121.920 0.000 125.460 1.120 ;
  LAYER ME2 ;
  RECT 121.920 0.000 125.460 1.120 ;
  LAYER ME1 ;
  RECT 121.920 0.000 125.460 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 100.220 0.000 103.760 1.120 ;
  LAYER ME3 ;
  RECT 100.220 0.000 103.760 1.120 ;
  LAYER ME2 ;
  RECT 100.220 0.000 103.760 1.120 ;
  LAYER ME1 ;
  RECT 100.220 0.000 103.760 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 83.480 0.000 87.020 1.120 ;
  LAYER ME3 ;
  RECT 83.480 0.000 87.020 1.120 ;
  LAYER ME2 ;
  RECT 83.480 0.000 87.020 1.120 ;
  LAYER ME1 ;
  RECT 83.480 0.000 87.020 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 56.820 0.000 60.360 1.120 ;
  LAYER ME3 ;
  RECT 56.820 0.000 60.360 1.120 ;
  LAYER ME2 ;
  RECT 56.820 0.000 60.360 1.120 ;
  LAYER ME1 ;
  RECT 56.820 0.000 60.360 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 35.740 0.000 39.280 1.120 ;
  LAYER ME3 ;
  RECT 35.740 0.000 39.280 1.120 ;
  LAYER ME2 ;
  RECT 35.740 0.000 39.280 1.120 ;
  LAYER ME1 ;
  RECT 35.740 0.000 39.280 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 14.040 0.000 17.580 1.120 ;
  LAYER ME3 ;
  RECT 14.040 0.000 17.580 1.120 ;
  LAYER ME2 ;
  RECT 14.040 0.000 17.580 1.120 ;
  LAYER ME1 ;
  RECT 14.040 0.000 17.580 1.120 ;
 END
END VCC
PIN DO15
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 292.080 0.000 293.200 1.120 ;
  LAYER ME3 ;
  RECT 292.080 0.000 293.200 1.120 ;
  LAYER ME2 ;
  RECT 292.080 0.000 293.200 1.120 ;
  LAYER ME1 ;
  RECT 292.080 0.000 293.200 1.120 ;
 END
END DO15
PIN DI15
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 284.020 0.000 285.140 1.120 ;
  LAYER ME3 ;
  RECT 284.020 0.000 285.140 1.120 ;
  LAYER ME2 ;
  RECT 284.020 0.000 285.140 1.120 ;
  LAYER ME1 ;
  RECT 284.020 0.000 285.140 1.120 ;
 END
END DI15
PIN DO14
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 279.060 0.000 280.180 1.120 ;
  LAYER ME3 ;
  RECT 279.060 0.000 280.180 1.120 ;
  LAYER ME2 ;
  RECT 279.060 0.000 280.180 1.120 ;
  LAYER ME1 ;
  RECT 279.060 0.000 280.180 1.120 ;
 END
END DO14
PIN DI14
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 270.380 0.000 271.500 1.120 ;
  LAYER ME3 ;
  RECT 270.380 0.000 271.500 1.120 ;
  LAYER ME2 ;
  RECT 270.380 0.000 271.500 1.120 ;
  LAYER ME1 ;
  RECT 270.380 0.000 271.500 1.120 ;
 END
END DI14
PIN DO13
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 262.320 0.000 263.440 1.120 ;
  LAYER ME3 ;
  RECT 262.320 0.000 263.440 1.120 ;
  LAYER ME2 ;
  RECT 262.320 0.000 263.440 1.120 ;
  LAYER ME1 ;
  RECT 262.320 0.000 263.440 1.120 ;
 END
END DO13
PIN DI13
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 253.640 0.000 254.760 1.120 ;
  LAYER ME3 ;
  RECT 253.640 0.000 254.760 1.120 ;
  LAYER ME2 ;
  RECT 253.640 0.000 254.760 1.120 ;
  LAYER ME1 ;
  RECT 253.640 0.000 254.760 1.120 ;
 END
END DI13
PIN DO12
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 248.680 0.000 249.800 1.120 ;
  LAYER ME3 ;
  RECT 248.680 0.000 249.800 1.120 ;
  LAYER ME2 ;
  RECT 248.680 0.000 249.800 1.120 ;
  LAYER ME1 ;
  RECT 248.680 0.000 249.800 1.120 ;
 END
END DO12
PIN DI12
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 240.620 0.000 241.740 1.120 ;
  LAYER ME3 ;
  RECT 240.620 0.000 241.740 1.120 ;
  LAYER ME2 ;
  RECT 240.620 0.000 241.740 1.120 ;
  LAYER ME1 ;
  RECT 240.620 0.000 241.740 1.120 ;
 END
END DI12
PIN DO11
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 235.660 0.000 236.780 1.120 ;
  LAYER ME3 ;
  RECT 235.660 0.000 236.780 1.120 ;
  LAYER ME2 ;
  RECT 235.660 0.000 236.780 1.120 ;
  LAYER ME1 ;
  RECT 235.660 0.000 236.780 1.120 ;
 END
END DO11
PIN DI11
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 226.980 0.000 228.100 1.120 ;
  LAYER ME3 ;
  RECT 226.980 0.000 228.100 1.120 ;
  LAYER ME2 ;
  RECT 226.980 0.000 228.100 1.120 ;
  LAYER ME1 ;
  RECT 226.980 0.000 228.100 1.120 ;
 END
END DI11
PIN DO10
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 222.020 0.000 223.140 1.120 ;
  LAYER ME3 ;
  RECT 222.020 0.000 223.140 1.120 ;
  LAYER ME2 ;
  RECT 222.020 0.000 223.140 1.120 ;
  LAYER ME1 ;
  RECT 222.020 0.000 223.140 1.120 ;
 END
END DO10
PIN DI10
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 213.960 0.000 215.080 1.120 ;
  LAYER ME3 ;
  RECT 213.960 0.000 215.080 1.120 ;
  LAYER ME2 ;
  RECT 213.960 0.000 215.080 1.120 ;
  LAYER ME1 ;
  RECT 213.960 0.000 215.080 1.120 ;
 END
END DI10
PIN DO9
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 205.900 0.000 207.020 1.120 ;
  LAYER ME3 ;
  RECT 205.900 0.000 207.020 1.120 ;
  LAYER ME2 ;
  RECT 205.900 0.000 207.020 1.120 ;
  LAYER ME1 ;
  RECT 205.900 0.000 207.020 1.120 ;
 END
END DO9
PIN DI9
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 197.220 0.000 198.340 1.120 ;
  LAYER ME3 ;
  RECT 197.220 0.000 198.340 1.120 ;
  LAYER ME2 ;
  RECT 197.220 0.000 198.340 1.120 ;
  LAYER ME1 ;
  RECT 197.220 0.000 198.340 1.120 ;
 END
END DI9
PIN DO8
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 192.260 0.000 193.380 1.120 ;
  LAYER ME3 ;
  RECT 192.260 0.000 193.380 1.120 ;
  LAYER ME2 ;
  RECT 192.260 0.000 193.380 1.120 ;
  LAYER ME1 ;
  RECT 192.260 0.000 193.380 1.120 ;
 END
END DO8
PIN DI8
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 184.200 0.000 185.320 1.120 ;
  LAYER ME3 ;
  RECT 184.200 0.000 185.320 1.120 ;
  LAYER ME2 ;
  RECT 184.200 0.000 185.320 1.120 ;
  LAYER ME1 ;
  RECT 184.200 0.000 185.320 1.120 ;
 END
END DI8
PIN A1
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 178.620 0.000 179.740 1.120 ;
  LAYER ME3 ;
  RECT 178.620 0.000 179.740 1.120 ;
  LAYER ME2 ;
  RECT 178.620 0.000 179.740 1.120 ;
  LAYER ME1 ;
  RECT 178.620 0.000 179.740 1.120 ;
 END
END A1
PIN WEB
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER ME4 ;
  RECT 176.760 0.000 177.880 1.120 ;
  LAYER ME3 ;
  RECT 176.760 0.000 177.880 1.120 ;
  LAYER ME2 ;
  RECT 176.760 0.000 177.880 1.120 ;
  LAYER ME1 ;
  RECT 176.760 0.000 177.880 1.120 ;
 END
END WEB
PIN OE
  DIRECTION INPUT ;
  CAPACITANCE 0.033 ;
 PORT
  LAYER ME4 ;
  RECT 171.800 0.000 172.920 1.120 ;
  LAYER ME3 ;
  RECT 171.800 0.000 172.920 1.120 ;
  LAYER ME2 ;
  RECT 171.800 0.000 172.920 1.120 ;
  LAYER ME1 ;
  RECT 171.800 0.000 172.920 1.120 ;
 END
END OE
PIN CS
  DIRECTION INPUT ;
  CAPACITANCE 0.123 ;
 PORT
  LAYER ME4 ;
  RECT 169.940 0.000 171.060 1.120 ;
  LAYER ME3 ;
  RECT 169.940 0.000 171.060 1.120 ;
  LAYER ME2 ;
  RECT 169.940 0.000 171.060 1.120 ;
  LAYER ME1 ;
  RECT 169.940 0.000 171.060 1.120 ;
 END
END CS
PIN A2
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 148.240 0.000 149.360 1.120 ;
  LAYER ME3 ;
  RECT 148.240 0.000 149.360 1.120 ;
  LAYER ME2 ;
  RECT 148.240 0.000 149.360 1.120 ;
  LAYER ME1 ;
  RECT 148.240 0.000 149.360 1.120 ;
 END
END A2
PIN CK
  DIRECTION INPUT ;
  CAPACITANCE 0.063 ;
 PORT
  LAYER ME4 ;
  RECT 145.140 0.000 146.260 1.120 ;
  LAYER ME3 ;
  RECT 145.140 0.000 146.260 1.120 ;
  LAYER ME2 ;
  RECT 145.140 0.000 146.260 1.120 ;
  LAYER ME1 ;
  RECT 145.140 0.000 146.260 1.120 ;
 END
END CK
PIN A0
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 142.660 0.000 143.780 1.120 ;
  LAYER ME3 ;
  RECT 142.660 0.000 143.780 1.120 ;
  LAYER ME2 ;
  RECT 142.660 0.000 143.780 1.120 ;
  LAYER ME1 ;
  RECT 142.660 0.000 143.780 1.120 ;
 END
END A0
PIN A3
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 138.320 0.000 139.440 1.120 ;
  LAYER ME3 ;
  RECT 138.320 0.000 139.440 1.120 ;
  LAYER ME2 ;
  RECT 138.320 0.000 139.440 1.120 ;
  LAYER ME1 ;
  RECT 138.320 0.000 139.440 1.120 ;
 END
END A3
PIN A4
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 130.880 0.000 132.000 1.120 ;
  LAYER ME3 ;
  RECT 130.880 0.000 132.000 1.120 ;
  LAYER ME2 ;
  RECT 130.880 0.000 132.000 1.120 ;
  LAYER ME1 ;
  RECT 130.880 0.000 132.000 1.120 ;
 END
END A4
PIN A5
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 127.780 0.000 128.900 1.120 ;
  LAYER ME3 ;
  RECT 127.780 0.000 128.900 1.120 ;
  LAYER ME2 ;
  RECT 127.780 0.000 128.900 1.120 ;
  LAYER ME1 ;
  RECT 127.780 0.000 128.900 1.120 ;
 END
END A5
PIN DO7
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 119.720 0.000 120.840 1.120 ;
  LAYER ME3 ;
  RECT 119.720 0.000 120.840 1.120 ;
  LAYER ME2 ;
  RECT 119.720 0.000 120.840 1.120 ;
  LAYER ME1 ;
  RECT 119.720 0.000 120.840 1.120 ;
 END
END DO7
PIN DI7
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 111.660 0.000 112.780 1.120 ;
  LAYER ME3 ;
  RECT 111.660 0.000 112.780 1.120 ;
  LAYER ME2 ;
  RECT 111.660 0.000 112.780 1.120 ;
  LAYER ME1 ;
  RECT 111.660 0.000 112.780 1.120 ;
 END
END DI7
PIN DO6
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 106.700 0.000 107.820 1.120 ;
  LAYER ME3 ;
  RECT 106.700 0.000 107.820 1.120 ;
  LAYER ME2 ;
  RECT 106.700 0.000 107.820 1.120 ;
  LAYER ME1 ;
  RECT 106.700 0.000 107.820 1.120 ;
 END
END DO6
PIN DI6
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 98.020 0.000 99.140 1.120 ;
  LAYER ME3 ;
  RECT 98.020 0.000 99.140 1.120 ;
  LAYER ME2 ;
  RECT 98.020 0.000 99.140 1.120 ;
  LAYER ME1 ;
  RECT 98.020 0.000 99.140 1.120 ;
 END
END DI6
PIN DO5
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 89.960 0.000 91.080 1.120 ;
  LAYER ME3 ;
  RECT 89.960 0.000 91.080 1.120 ;
  LAYER ME2 ;
  RECT 89.960 0.000 91.080 1.120 ;
  LAYER ME1 ;
  RECT 89.960 0.000 91.080 1.120 ;
 END
END DO5
PIN DI5
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 81.280 0.000 82.400 1.120 ;
  LAYER ME3 ;
  RECT 81.280 0.000 82.400 1.120 ;
  LAYER ME2 ;
  RECT 81.280 0.000 82.400 1.120 ;
  LAYER ME1 ;
  RECT 81.280 0.000 82.400 1.120 ;
 END
END DI5
PIN DO4
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 76.320 0.000 77.440 1.120 ;
  LAYER ME3 ;
  RECT 76.320 0.000 77.440 1.120 ;
  LAYER ME2 ;
  RECT 76.320 0.000 77.440 1.120 ;
  LAYER ME1 ;
  RECT 76.320 0.000 77.440 1.120 ;
 END
END DO4
PIN DI4
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 68.260 0.000 69.380 1.120 ;
  LAYER ME3 ;
  RECT 68.260 0.000 69.380 1.120 ;
  LAYER ME2 ;
  RECT 68.260 0.000 69.380 1.120 ;
  LAYER ME1 ;
  RECT 68.260 0.000 69.380 1.120 ;
 END
END DI4
PIN DO3
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 63.300 0.000 64.420 1.120 ;
  LAYER ME3 ;
  RECT 63.300 0.000 64.420 1.120 ;
  LAYER ME2 ;
  RECT 63.300 0.000 64.420 1.120 ;
  LAYER ME1 ;
  RECT 63.300 0.000 64.420 1.120 ;
 END
END DO3
PIN DI3
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 54.620 0.000 55.740 1.120 ;
  LAYER ME3 ;
  RECT 54.620 0.000 55.740 1.120 ;
  LAYER ME2 ;
  RECT 54.620 0.000 55.740 1.120 ;
  LAYER ME1 ;
  RECT 54.620 0.000 55.740 1.120 ;
 END
END DI3
PIN DO2
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 50.280 0.000 51.400 1.120 ;
  LAYER ME3 ;
  RECT 50.280 0.000 51.400 1.120 ;
  LAYER ME2 ;
  RECT 50.280 0.000 51.400 1.120 ;
  LAYER ME1 ;
  RECT 50.280 0.000 51.400 1.120 ;
 END
END DO2
PIN DI2
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 41.600 0.000 42.720 1.120 ;
  LAYER ME3 ;
  RECT 41.600 0.000 42.720 1.120 ;
  LAYER ME2 ;
  RECT 41.600 0.000 42.720 1.120 ;
  LAYER ME1 ;
  RECT 41.600 0.000 42.720 1.120 ;
 END
END DI2
PIN DO1
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 33.540 0.000 34.660 1.120 ;
  LAYER ME3 ;
  RECT 33.540 0.000 34.660 1.120 ;
  LAYER ME2 ;
  RECT 33.540 0.000 34.660 1.120 ;
  LAYER ME1 ;
  RECT 33.540 0.000 34.660 1.120 ;
 END
END DO1
PIN DI1
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 24.860 0.000 25.980 1.120 ;
  LAYER ME3 ;
  RECT 24.860 0.000 25.980 1.120 ;
  LAYER ME2 ;
  RECT 24.860 0.000 25.980 1.120 ;
  LAYER ME1 ;
  RECT 24.860 0.000 25.980 1.120 ;
 END
END DI1
PIN DO0
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 19.900 0.000 21.020 1.120 ;
  LAYER ME3 ;
  RECT 19.900 0.000 21.020 1.120 ;
  LAYER ME2 ;
  RECT 19.900 0.000 21.020 1.120 ;
  LAYER ME1 ;
  RECT 19.900 0.000 21.020 1.120 ;
 END
END DO0
PIN DI0
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 11.840 0.000 12.960 1.120 ;
  LAYER ME3 ;
  RECT 11.840 0.000 12.960 1.120 ;
  LAYER ME2 ;
  RECT 11.840 0.000 12.960 1.120 ;
  LAYER ME1 ;
  RECT 11.840 0.000 12.960 1.120 ;
 END
END DI0
OBS
  LAYER ME1 SPACING 0.280 ;
  RECT 0.000 0.140 305.660 156.800 ;
  LAYER ME2 SPACING 0.320 ;
  RECT 0.000 0.140 305.660 156.800 ;
  LAYER ME3 SPACING 0.320 ;
  RECT 0.000 0.140 305.660 156.800 ;
  LAYER ME4 SPACING 0.600 ;
  RECT 0.000 0.140 305.660 156.800 ;
  LAYER VI1 ;
  RECT 0.000 0.140 305.660 156.800 ;
  LAYER VI2 ;
  RECT 0.000 0.140 305.660 156.800 ;
  LAYER VI3 ;
  RECT 0.000 0.140 305.660 156.800 ;
END
END Memory_16_64
END LIBRARY



